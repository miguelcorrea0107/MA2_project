magic
tech sky130A
magscale 1 2
timestamp 1716644424
<< metal3 >>
rect -2786 2592 2786 2640
rect -2786 2528 2702 2592
rect 2766 2528 2786 2592
rect -2786 2512 2786 2528
rect -2786 2448 2702 2512
rect 2766 2448 2786 2512
rect -2786 2432 2786 2448
rect -2786 2368 2702 2432
rect 2766 2368 2786 2432
rect -2786 2352 2786 2368
rect -2786 2288 2702 2352
rect 2766 2288 2786 2352
rect -2786 2272 2786 2288
rect -2786 2208 2702 2272
rect 2766 2208 2786 2272
rect -2786 2192 2786 2208
rect -2786 2128 2702 2192
rect 2766 2128 2786 2192
rect -2786 2112 2786 2128
rect -2786 2048 2702 2112
rect 2766 2048 2786 2112
rect -2786 2032 2786 2048
rect -2786 1968 2702 2032
rect 2766 1968 2786 2032
rect -2786 1952 2786 1968
rect -2786 1888 2702 1952
rect 2766 1888 2786 1952
rect -2786 1872 2786 1888
rect -2786 1808 2702 1872
rect 2766 1808 2786 1872
rect -2786 1792 2786 1808
rect -2786 1728 2702 1792
rect 2766 1728 2786 1792
rect -2786 1712 2786 1728
rect -2786 1648 2702 1712
rect 2766 1648 2786 1712
rect -2786 1632 2786 1648
rect -2786 1568 2702 1632
rect 2766 1568 2786 1632
rect -2786 1552 2786 1568
rect -2786 1488 2702 1552
rect 2766 1488 2786 1552
rect -2786 1472 2786 1488
rect -2786 1408 2702 1472
rect 2766 1408 2786 1472
rect -2786 1392 2786 1408
rect -2786 1328 2702 1392
rect 2766 1328 2786 1392
rect -2786 1312 2786 1328
rect -2786 1248 2702 1312
rect 2766 1248 2786 1312
rect -2786 1232 2786 1248
rect -2786 1168 2702 1232
rect 2766 1168 2786 1232
rect -2786 1152 2786 1168
rect -2786 1088 2702 1152
rect 2766 1088 2786 1152
rect -2786 1072 2786 1088
rect -2786 1008 2702 1072
rect 2766 1008 2786 1072
rect -2786 992 2786 1008
rect -2786 928 2702 992
rect 2766 928 2786 992
rect -2786 912 2786 928
rect -2786 848 2702 912
rect 2766 848 2786 912
rect -2786 832 2786 848
rect -2786 768 2702 832
rect 2766 768 2786 832
rect -2786 752 2786 768
rect -2786 688 2702 752
rect 2766 688 2786 752
rect -2786 672 2786 688
rect -2786 608 2702 672
rect 2766 608 2786 672
rect -2786 592 2786 608
rect -2786 528 2702 592
rect 2766 528 2786 592
rect -2786 512 2786 528
rect -2786 448 2702 512
rect 2766 448 2786 512
rect -2786 432 2786 448
rect -2786 368 2702 432
rect 2766 368 2786 432
rect -2786 352 2786 368
rect -2786 288 2702 352
rect 2766 288 2786 352
rect -2786 272 2786 288
rect -2786 208 2702 272
rect 2766 208 2786 272
rect -2786 192 2786 208
rect -2786 128 2702 192
rect 2766 128 2786 192
rect -2786 112 2786 128
rect -2786 48 2702 112
rect 2766 48 2786 112
rect -2786 32 2786 48
rect -2786 -32 2702 32
rect 2766 -32 2786 32
rect -2786 -48 2786 -32
rect -2786 -112 2702 -48
rect 2766 -112 2786 -48
rect -2786 -128 2786 -112
rect -2786 -192 2702 -128
rect 2766 -192 2786 -128
rect -2786 -208 2786 -192
rect -2786 -272 2702 -208
rect 2766 -272 2786 -208
rect -2786 -288 2786 -272
rect -2786 -352 2702 -288
rect 2766 -352 2786 -288
rect -2786 -368 2786 -352
rect -2786 -432 2702 -368
rect 2766 -432 2786 -368
rect -2786 -448 2786 -432
rect -2786 -512 2702 -448
rect 2766 -512 2786 -448
rect -2786 -528 2786 -512
rect -2786 -592 2702 -528
rect 2766 -592 2786 -528
rect -2786 -608 2786 -592
rect -2786 -672 2702 -608
rect 2766 -672 2786 -608
rect -2786 -688 2786 -672
rect -2786 -752 2702 -688
rect 2766 -752 2786 -688
rect -2786 -768 2786 -752
rect -2786 -832 2702 -768
rect 2766 -832 2786 -768
rect -2786 -848 2786 -832
rect -2786 -912 2702 -848
rect 2766 -912 2786 -848
rect -2786 -928 2786 -912
rect -2786 -992 2702 -928
rect 2766 -992 2786 -928
rect -2786 -1008 2786 -992
rect -2786 -1072 2702 -1008
rect 2766 -1072 2786 -1008
rect -2786 -1088 2786 -1072
rect -2786 -1152 2702 -1088
rect 2766 -1152 2786 -1088
rect -2786 -1168 2786 -1152
rect -2786 -1232 2702 -1168
rect 2766 -1232 2786 -1168
rect -2786 -1248 2786 -1232
rect -2786 -1312 2702 -1248
rect 2766 -1312 2786 -1248
rect -2786 -1328 2786 -1312
rect -2786 -1392 2702 -1328
rect 2766 -1392 2786 -1328
rect -2786 -1408 2786 -1392
rect -2786 -1472 2702 -1408
rect 2766 -1472 2786 -1408
rect -2786 -1488 2786 -1472
rect -2786 -1552 2702 -1488
rect 2766 -1552 2786 -1488
rect -2786 -1568 2786 -1552
rect -2786 -1632 2702 -1568
rect 2766 -1632 2786 -1568
rect -2786 -1648 2786 -1632
rect -2786 -1712 2702 -1648
rect 2766 -1712 2786 -1648
rect -2786 -1728 2786 -1712
rect -2786 -1792 2702 -1728
rect 2766 -1792 2786 -1728
rect -2786 -1808 2786 -1792
rect -2786 -1872 2702 -1808
rect 2766 -1872 2786 -1808
rect -2786 -1888 2786 -1872
rect -2786 -1952 2702 -1888
rect 2766 -1952 2786 -1888
rect -2786 -1968 2786 -1952
rect -2786 -2032 2702 -1968
rect 2766 -2032 2786 -1968
rect -2786 -2048 2786 -2032
rect -2786 -2112 2702 -2048
rect 2766 -2112 2786 -2048
rect -2786 -2128 2786 -2112
rect -2786 -2192 2702 -2128
rect 2766 -2192 2786 -2128
rect -2786 -2208 2786 -2192
rect -2786 -2272 2702 -2208
rect 2766 -2272 2786 -2208
rect -2786 -2288 2786 -2272
rect -2786 -2352 2702 -2288
rect 2766 -2352 2786 -2288
rect -2786 -2368 2786 -2352
rect -2786 -2432 2702 -2368
rect 2766 -2432 2786 -2368
rect -2786 -2448 2786 -2432
rect -2786 -2512 2702 -2448
rect 2766 -2512 2786 -2448
rect -2786 -2528 2786 -2512
rect -2786 -2592 2702 -2528
rect 2766 -2592 2786 -2528
rect -2786 -2640 2786 -2592
<< via3 >>
rect 2702 2528 2766 2592
rect 2702 2448 2766 2512
rect 2702 2368 2766 2432
rect 2702 2288 2766 2352
rect 2702 2208 2766 2272
rect 2702 2128 2766 2192
rect 2702 2048 2766 2112
rect 2702 1968 2766 2032
rect 2702 1888 2766 1952
rect 2702 1808 2766 1872
rect 2702 1728 2766 1792
rect 2702 1648 2766 1712
rect 2702 1568 2766 1632
rect 2702 1488 2766 1552
rect 2702 1408 2766 1472
rect 2702 1328 2766 1392
rect 2702 1248 2766 1312
rect 2702 1168 2766 1232
rect 2702 1088 2766 1152
rect 2702 1008 2766 1072
rect 2702 928 2766 992
rect 2702 848 2766 912
rect 2702 768 2766 832
rect 2702 688 2766 752
rect 2702 608 2766 672
rect 2702 528 2766 592
rect 2702 448 2766 512
rect 2702 368 2766 432
rect 2702 288 2766 352
rect 2702 208 2766 272
rect 2702 128 2766 192
rect 2702 48 2766 112
rect 2702 -32 2766 32
rect 2702 -112 2766 -48
rect 2702 -192 2766 -128
rect 2702 -272 2766 -208
rect 2702 -352 2766 -288
rect 2702 -432 2766 -368
rect 2702 -512 2766 -448
rect 2702 -592 2766 -528
rect 2702 -672 2766 -608
rect 2702 -752 2766 -688
rect 2702 -832 2766 -768
rect 2702 -912 2766 -848
rect 2702 -992 2766 -928
rect 2702 -1072 2766 -1008
rect 2702 -1152 2766 -1088
rect 2702 -1232 2766 -1168
rect 2702 -1312 2766 -1248
rect 2702 -1392 2766 -1328
rect 2702 -1472 2766 -1408
rect 2702 -1552 2766 -1488
rect 2702 -1632 2766 -1568
rect 2702 -1712 2766 -1648
rect 2702 -1792 2766 -1728
rect 2702 -1872 2766 -1808
rect 2702 -1952 2766 -1888
rect 2702 -2032 2766 -1968
rect 2702 -2112 2766 -2048
rect 2702 -2192 2766 -2128
rect 2702 -2272 2766 -2208
rect 2702 -2352 2766 -2288
rect 2702 -2432 2766 -2368
rect 2702 -2512 2766 -2448
rect 2702 -2592 2766 -2528
<< mimcap >>
rect -2746 2552 2454 2600
rect -2746 -2552 -2698 2552
rect 2406 -2552 2454 2552
rect -2746 -2600 2454 -2552
<< mimcapcontact >>
rect -2698 -2552 2406 2552
<< metal4 >>
rect 2686 2592 2782 2628
rect -2707 2552 2415 2561
rect -2707 -2552 -2698 2552
rect 2406 -2552 2415 2552
rect -2707 -2561 2415 -2552
rect 2686 2528 2702 2592
rect 2766 2528 2782 2592
rect 2686 2512 2782 2528
rect 2686 2448 2702 2512
rect 2766 2448 2782 2512
rect 2686 2432 2782 2448
rect 2686 2368 2702 2432
rect 2766 2368 2782 2432
rect 2686 2352 2782 2368
rect 2686 2288 2702 2352
rect 2766 2288 2782 2352
rect 2686 2272 2782 2288
rect 2686 2208 2702 2272
rect 2766 2208 2782 2272
rect 2686 2192 2782 2208
rect 2686 2128 2702 2192
rect 2766 2128 2782 2192
rect 2686 2112 2782 2128
rect 2686 2048 2702 2112
rect 2766 2048 2782 2112
rect 2686 2032 2782 2048
rect 2686 1968 2702 2032
rect 2766 1968 2782 2032
rect 2686 1952 2782 1968
rect 2686 1888 2702 1952
rect 2766 1888 2782 1952
rect 2686 1872 2782 1888
rect 2686 1808 2702 1872
rect 2766 1808 2782 1872
rect 2686 1792 2782 1808
rect 2686 1728 2702 1792
rect 2766 1728 2782 1792
rect 2686 1712 2782 1728
rect 2686 1648 2702 1712
rect 2766 1648 2782 1712
rect 2686 1632 2782 1648
rect 2686 1568 2702 1632
rect 2766 1568 2782 1632
rect 2686 1552 2782 1568
rect 2686 1488 2702 1552
rect 2766 1488 2782 1552
rect 2686 1472 2782 1488
rect 2686 1408 2702 1472
rect 2766 1408 2782 1472
rect 2686 1392 2782 1408
rect 2686 1328 2702 1392
rect 2766 1328 2782 1392
rect 2686 1312 2782 1328
rect 2686 1248 2702 1312
rect 2766 1248 2782 1312
rect 2686 1232 2782 1248
rect 2686 1168 2702 1232
rect 2766 1168 2782 1232
rect 2686 1152 2782 1168
rect 2686 1088 2702 1152
rect 2766 1088 2782 1152
rect 2686 1072 2782 1088
rect 2686 1008 2702 1072
rect 2766 1008 2782 1072
rect 2686 992 2782 1008
rect 2686 928 2702 992
rect 2766 928 2782 992
rect 2686 912 2782 928
rect 2686 848 2702 912
rect 2766 848 2782 912
rect 2686 832 2782 848
rect 2686 768 2702 832
rect 2766 768 2782 832
rect 2686 752 2782 768
rect 2686 688 2702 752
rect 2766 688 2782 752
rect 2686 672 2782 688
rect 2686 608 2702 672
rect 2766 608 2782 672
rect 2686 592 2782 608
rect 2686 528 2702 592
rect 2766 528 2782 592
rect 2686 512 2782 528
rect 2686 448 2702 512
rect 2766 448 2782 512
rect 2686 432 2782 448
rect 2686 368 2702 432
rect 2766 368 2782 432
rect 2686 352 2782 368
rect 2686 288 2702 352
rect 2766 288 2782 352
rect 2686 272 2782 288
rect 2686 208 2702 272
rect 2766 208 2782 272
rect 2686 192 2782 208
rect 2686 128 2702 192
rect 2766 128 2782 192
rect 2686 112 2782 128
rect 2686 48 2702 112
rect 2766 48 2782 112
rect 2686 32 2782 48
rect 2686 -32 2702 32
rect 2766 -32 2782 32
rect 2686 -48 2782 -32
rect 2686 -112 2702 -48
rect 2766 -112 2782 -48
rect 2686 -128 2782 -112
rect 2686 -192 2702 -128
rect 2766 -192 2782 -128
rect 2686 -208 2782 -192
rect 2686 -272 2702 -208
rect 2766 -272 2782 -208
rect 2686 -288 2782 -272
rect 2686 -352 2702 -288
rect 2766 -352 2782 -288
rect 2686 -368 2782 -352
rect 2686 -432 2702 -368
rect 2766 -432 2782 -368
rect 2686 -448 2782 -432
rect 2686 -512 2702 -448
rect 2766 -512 2782 -448
rect 2686 -528 2782 -512
rect 2686 -592 2702 -528
rect 2766 -592 2782 -528
rect 2686 -608 2782 -592
rect 2686 -672 2702 -608
rect 2766 -672 2782 -608
rect 2686 -688 2782 -672
rect 2686 -752 2702 -688
rect 2766 -752 2782 -688
rect 2686 -768 2782 -752
rect 2686 -832 2702 -768
rect 2766 -832 2782 -768
rect 2686 -848 2782 -832
rect 2686 -912 2702 -848
rect 2766 -912 2782 -848
rect 2686 -928 2782 -912
rect 2686 -992 2702 -928
rect 2766 -992 2782 -928
rect 2686 -1008 2782 -992
rect 2686 -1072 2702 -1008
rect 2766 -1072 2782 -1008
rect 2686 -1088 2782 -1072
rect 2686 -1152 2702 -1088
rect 2766 -1152 2782 -1088
rect 2686 -1168 2782 -1152
rect 2686 -1232 2702 -1168
rect 2766 -1232 2782 -1168
rect 2686 -1248 2782 -1232
rect 2686 -1312 2702 -1248
rect 2766 -1312 2782 -1248
rect 2686 -1328 2782 -1312
rect 2686 -1392 2702 -1328
rect 2766 -1392 2782 -1328
rect 2686 -1408 2782 -1392
rect 2686 -1472 2702 -1408
rect 2766 -1472 2782 -1408
rect 2686 -1488 2782 -1472
rect 2686 -1552 2702 -1488
rect 2766 -1552 2782 -1488
rect 2686 -1568 2782 -1552
rect 2686 -1632 2702 -1568
rect 2766 -1632 2782 -1568
rect 2686 -1648 2782 -1632
rect 2686 -1712 2702 -1648
rect 2766 -1712 2782 -1648
rect 2686 -1728 2782 -1712
rect 2686 -1792 2702 -1728
rect 2766 -1792 2782 -1728
rect 2686 -1808 2782 -1792
rect 2686 -1872 2702 -1808
rect 2766 -1872 2782 -1808
rect 2686 -1888 2782 -1872
rect 2686 -1952 2702 -1888
rect 2766 -1952 2782 -1888
rect 2686 -1968 2782 -1952
rect 2686 -2032 2702 -1968
rect 2766 -2032 2782 -1968
rect 2686 -2048 2782 -2032
rect 2686 -2112 2702 -2048
rect 2766 -2112 2782 -2048
rect 2686 -2128 2782 -2112
rect 2686 -2192 2702 -2128
rect 2766 -2192 2782 -2128
rect 2686 -2208 2782 -2192
rect 2686 -2272 2702 -2208
rect 2766 -2272 2782 -2208
rect 2686 -2288 2782 -2272
rect 2686 -2352 2702 -2288
rect 2766 -2352 2782 -2288
rect 2686 -2368 2782 -2352
rect 2686 -2432 2702 -2368
rect 2766 -2432 2782 -2368
rect 2686 -2448 2782 -2432
rect 2686 -2512 2702 -2448
rect 2766 -2512 2782 -2448
rect 2686 -2528 2782 -2512
rect 2686 -2592 2702 -2528
rect 2766 -2592 2782 -2528
rect 2686 -2628 2782 -2592
<< properties >>
string FIXED_BBOX -2786 -2640 2494 2640
<< end >>
