magic
tech sky130A
magscale 1 2
timestamp 1716644424
<< error_p >>
rect -299 2581 -241 2587
rect -83 2581 -25 2587
rect 133 2581 191 2587
rect 349 2581 407 2587
rect -299 2547 -287 2581
rect -83 2547 -71 2581
rect 133 2547 145 2581
rect 349 2547 361 2581
rect -299 2541 -241 2547
rect -83 2541 -25 2547
rect 133 2541 191 2547
rect 349 2541 407 2547
rect -407 -2547 -349 -2541
rect -191 -2547 -133 -2541
rect 25 -2547 83 -2541
rect 241 -2547 299 -2541
rect -407 -2581 -395 -2547
rect -191 -2581 -179 -2547
rect 25 -2581 37 -2547
rect 241 -2581 253 -2547
rect -407 -2587 -349 -2581
rect -191 -2587 -133 -2581
rect 25 -2587 83 -2581
rect 241 -2587 299 -2581
<< nwell >>
rect -599 -2719 599 2719
<< pmos >>
rect -403 -2500 -353 2500
rect -295 -2500 -245 2500
rect -187 -2500 -137 2500
rect -79 -2500 -29 2500
rect 29 -2500 79 2500
rect 137 -2500 187 2500
rect 245 -2500 295 2500
rect 353 -2500 403 2500
<< pdiff >>
rect -461 2465 -403 2500
rect -461 2431 -449 2465
rect -415 2431 -403 2465
rect -461 2397 -403 2431
rect -461 2363 -449 2397
rect -415 2363 -403 2397
rect -461 2329 -403 2363
rect -461 2295 -449 2329
rect -415 2295 -403 2329
rect -461 2261 -403 2295
rect -461 2227 -449 2261
rect -415 2227 -403 2261
rect -461 2193 -403 2227
rect -461 2159 -449 2193
rect -415 2159 -403 2193
rect -461 2125 -403 2159
rect -461 2091 -449 2125
rect -415 2091 -403 2125
rect -461 2057 -403 2091
rect -461 2023 -449 2057
rect -415 2023 -403 2057
rect -461 1989 -403 2023
rect -461 1955 -449 1989
rect -415 1955 -403 1989
rect -461 1921 -403 1955
rect -461 1887 -449 1921
rect -415 1887 -403 1921
rect -461 1853 -403 1887
rect -461 1819 -449 1853
rect -415 1819 -403 1853
rect -461 1785 -403 1819
rect -461 1751 -449 1785
rect -415 1751 -403 1785
rect -461 1717 -403 1751
rect -461 1683 -449 1717
rect -415 1683 -403 1717
rect -461 1649 -403 1683
rect -461 1615 -449 1649
rect -415 1615 -403 1649
rect -461 1581 -403 1615
rect -461 1547 -449 1581
rect -415 1547 -403 1581
rect -461 1513 -403 1547
rect -461 1479 -449 1513
rect -415 1479 -403 1513
rect -461 1445 -403 1479
rect -461 1411 -449 1445
rect -415 1411 -403 1445
rect -461 1377 -403 1411
rect -461 1343 -449 1377
rect -415 1343 -403 1377
rect -461 1309 -403 1343
rect -461 1275 -449 1309
rect -415 1275 -403 1309
rect -461 1241 -403 1275
rect -461 1207 -449 1241
rect -415 1207 -403 1241
rect -461 1173 -403 1207
rect -461 1139 -449 1173
rect -415 1139 -403 1173
rect -461 1105 -403 1139
rect -461 1071 -449 1105
rect -415 1071 -403 1105
rect -461 1037 -403 1071
rect -461 1003 -449 1037
rect -415 1003 -403 1037
rect -461 969 -403 1003
rect -461 935 -449 969
rect -415 935 -403 969
rect -461 901 -403 935
rect -461 867 -449 901
rect -415 867 -403 901
rect -461 833 -403 867
rect -461 799 -449 833
rect -415 799 -403 833
rect -461 765 -403 799
rect -461 731 -449 765
rect -415 731 -403 765
rect -461 697 -403 731
rect -461 663 -449 697
rect -415 663 -403 697
rect -461 629 -403 663
rect -461 595 -449 629
rect -415 595 -403 629
rect -461 561 -403 595
rect -461 527 -449 561
rect -415 527 -403 561
rect -461 493 -403 527
rect -461 459 -449 493
rect -415 459 -403 493
rect -461 425 -403 459
rect -461 391 -449 425
rect -415 391 -403 425
rect -461 357 -403 391
rect -461 323 -449 357
rect -415 323 -403 357
rect -461 289 -403 323
rect -461 255 -449 289
rect -415 255 -403 289
rect -461 221 -403 255
rect -461 187 -449 221
rect -415 187 -403 221
rect -461 153 -403 187
rect -461 119 -449 153
rect -415 119 -403 153
rect -461 85 -403 119
rect -461 51 -449 85
rect -415 51 -403 85
rect -461 17 -403 51
rect -461 -17 -449 17
rect -415 -17 -403 17
rect -461 -51 -403 -17
rect -461 -85 -449 -51
rect -415 -85 -403 -51
rect -461 -119 -403 -85
rect -461 -153 -449 -119
rect -415 -153 -403 -119
rect -461 -187 -403 -153
rect -461 -221 -449 -187
rect -415 -221 -403 -187
rect -461 -255 -403 -221
rect -461 -289 -449 -255
rect -415 -289 -403 -255
rect -461 -323 -403 -289
rect -461 -357 -449 -323
rect -415 -357 -403 -323
rect -461 -391 -403 -357
rect -461 -425 -449 -391
rect -415 -425 -403 -391
rect -461 -459 -403 -425
rect -461 -493 -449 -459
rect -415 -493 -403 -459
rect -461 -527 -403 -493
rect -461 -561 -449 -527
rect -415 -561 -403 -527
rect -461 -595 -403 -561
rect -461 -629 -449 -595
rect -415 -629 -403 -595
rect -461 -663 -403 -629
rect -461 -697 -449 -663
rect -415 -697 -403 -663
rect -461 -731 -403 -697
rect -461 -765 -449 -731
rect -415 -765 -403 -731
rect -461 -799 -403 -765
rect -461 -833 -449 -799
rect -415 -833 -403 -799
rect -461 -867 -403 -833
rect -461 -901 -449 -867
rect -415 -901 -403 -867
rect -461 -935 -403 -901
rect -461 -969 -449 -935
rect -415 -969 -403 -935
rect -461 -1003 -403 -969
rect -461 -1037 -449 -1003
rect -415 -1037 -403 -1003
rect -461 -1071 -403 -1037
rect -461 -1105 -449 -1071
rect -415 -1105 -403 -1071
rect -461 -1139 -403 -1105
rect -461 -1173 -449 -1139
rect -415 -1173 -403 -1139
rect -461 -1207 -403 -1173
rect -461 -1241 -449 -1207
rect -415 -1241 -403 -1207
rect -461 -1275 -403 -1241
rect -461 -1309 -449 -1275
rect -415 -1309 -403 -1275
rect -461 -1343 -403 -1309
rect -461 -1377 -449 -1343
rect -415 -1377 -403 -1343
rect -461 -1411 -403 -1377
rect -461 -1445 -449 -1411
rect -415 -1445 -403 -1411
rect -461 -1479 -403 -1445
rect -461 -1513 -449 -1479
rect -415 -1513 -403 -1479
rect -461 -1547 -403 -1513
rect -461 -1581 -449 -1547
rect -415 -1581 -403 -1547
rect -461 -1615 -403 -1581
rect -461 -1649 -449 -1615
rect -415 -1649 -403 -1615
rect -461 -1683 -403 -1649
rect -461 -1717 -449 -1683
rect -415 -1717 -403 -1683
rect -461 -1751 -403 -1717
rect -461 -1785 -449 -1751
rect -415 -1785 -403 -1751
rect -461 -1819 -403 -1785
rect -461 -1853 -449 -1819
rect -415 -1853 -403 -1819
rect -461 -1887 -403 -1853
rect -461 -1921 -449 -1887
rect -415 -1921 -403 -1887
rect -461 -1955 -403 -1921
rect -461 -1989 -449 -1955
rect -415 -1989 -403 -1955
rect -461 -2023 -403 -1989
rect -461 -2057 -449 -2023
rect -415 -2057 -403 -2023
rect -461 -2091 -403 -2057
rect -461 -2125 -449 -2091
rect -415 -2125 -403 -2091
rect -461 -2159 -403 -2125
rect -461 -2193 -449 -2159
rect -415 -2193 -403 -2159
rect -461 -2227 -403 -2193
rect -461 -2261 -449 -2227
rect -415 -2261 -403 -2227
rect -461 -2295 -403 -2261
rect -461 -2329 -449 -2295
rect -415 -2329 -403 -2295
rect -461 -2363 -403 -2329
rect -461 -2397 -449 -2363
rect -415 -2397 -403 -2363
rect -461 -2431 -403 -2397
rect -461 -2465 -449 -2431
rect -415 -2465 -403 -2431
rect -461 -2500 -403 -2465
rect -353 2465 -295 2500
rect -353 2431 -341 2465
rect -307 2431 -295 2465
rect -353 2397 -295 2431
rect -353 2363 -341 2397
rect -307 2363 -295 2397
rect -353 2329 -295 2363
rect -353 2295 -341 2329
rect -307 2295 -295 2329
rect -353 2261 -295 2295
rect -353 2227 -341 2261
rect -307 2227 -295 2261
rect -353 2193 -295 2227
rect -353 2159 -341 2193
rect -307 2159 -295 2193
rect -353 2125 -295 2159
rect -353 2091 -341 2125
rect -307 2091 -295 2125
rect -353 2057 -295 2091
rect -353 2023 -341 2057
rect -307 2023 -295 2057
rect -353 1989 -295 2023
rect -353 1955 -341 1989
rect -307 1955 -295 1989
rect -353 1921 -295 1955
rect -353 1887 -341 1921
rect -307 1887 -295 1921
rect -353 1853 -295 1887
rect -353 1819 -341 1853
rect -307 1819 -295 1853
rect -353 1785 -295 1819
rect -353 1751 -341 1785
rect -307 1751 -295 1785
rect -353 1717 -295 1751
rect -353 1683 -341 1717
rect -307 1683 -295 1717
rect -353 1649 -295 1683
rect -353 1615 -341 1649
rect -307 1615 -295 1649
rect -353 1581 -295 1615
rect -353 1547 -341 1581
rect -307 1547 -295 1581
rect -353 1513 -295 1547
rect -353 1479 -341 1513
rect -307 1479 -295 1513
rect -353 1445 -295 1479
rect -353 1411 -341 1445
rect -307 1411 -295 1445
rect -353 1377 -295 1411
rect -353 1343 -341 1377
rect -307 1343 -295 1377
rect -353 1309 -295 1343
rect -353 1275 -341 1309
rect -307 1275 -295 1309
rect -353 1241 -295 1275
rect -353 1207 -341 1241
rect -307 1207 -295 1241
rect -353 1173 -295 1207
rect -353 1139 -341 1173
rect -307 1139 -295 1173
rect -353 1105 -295 1139
rect -353 1071 -341 1105
rect -307 1071 -295 1105
rect -353 1037 -295 1071
rect -353 1003 -341 1037
rect -307 1003 -295 1037
rect -353 969 -295 1003
rect -353 935 -341 969
rect -307 935 -295 969
rect -353 901 -295 935
rect -353 867 -341 901
rect -307 867 -295 901
rect -353 833 -295 867
rect -353 799 -341 833
rect -307 799 -295 833
rect -353 765 -295 799
rect -353 731 -341 765
rect -307 731 -295 765
rect -353 697 -295 731
rect -353 663 -341 697
rect -307 663 -295 697
rect -353 629 -295 663
rect -353 595 -341 629
rect -307 595 -295 629
rect -353 561 -295 595
rect -353 527 -341 561
rect -307 527 -295 561
rect -353 493 -295 527
rect -353 459 -341 493
rect -307 459 -295 493
rect -353 425 -295 459
rect -353 391 -341 425
rect -307 391 -295 425
rect -353 357 -295 391
rect -353 323 -341 357
rect -307 323 -295 357
rect -353 289 -295 323
rect -353 255 -341 289
rect -307 255 -295 289
rect -353 221 -295 255
rect -353 187 -341 221
rect -307 187 -295 221
rect -353 153 -295 187
rect -353 119 -341 153
rect -307 119 -295 153
rect -353 85 -295 119
rect -353 51 -341 85
rect -307 51 -295 85
rect -353 17 -295 51
rect -353 -17 -341 17
rect -307 -17 -295 17
rect -353 -51 -295 -17
rect -353 -85 -341 -51
rect -307 -85 -295 -51
rect -353 -119 -295 -85
rect -353 -153 -341 -119
rect -307 -153 -295 -119
rect -353 -187 -295 -153
rect -353 -221 -341 -187
rect -307 -221 -295 -187
rect -353 -255 -295 -221
rect -353 -289 -341 -255
rect -307 -289 -295 -255
rect -353 -323 -295 -289
rect -353 -357 -341 -323
rect -307 -357 -295 -323
rect -353 -391 -295 -357
rect -353 -425 -341 -391
rect -307 -425 -295 -391
rect -353 -459 -295 -425
rect -353 -493 -341 -459
rect -307 -493 -295 -459
rect -353 -527 -295 -493
rect -353 -561 -341 -527
rect -307 -561 -295 -527
rect -353 -595 -295 -561
rect -353 -629 -341 -595
rect -307 -629 -295 -595
rect -353 -663 -295 -629
rect -353 -697 -341 -663
rect -307 -697 -295 -663
rect -353 -731 -295 -697
rect -353 -765 -341 -731
rect -307 -765 -295 -731
rect -353 -799 -295 -765
rect -353 -833 -341 -799
rect -307 -833 -295 -799
rect -353 -867 -295 -833
rect -353 -901 -341 -867
rect -307 -901 -295 -867
rect -353 -935 -295 -901
rect -353 -969 -341 -935
rect -307 -969 -295 -935
rect -353 -1003 -295 -969
rect -353 -1037 -341 -1003
rect -307 -1037 -295 -1003
rect -353 -1071 -295 -1037
rect -353 -1105 -341 -1071
rect -307 -1105 -295 -1071
rect -353 -1139 -295 -1105
rect -353 -1173 -341 -1139
rect -307 -1173 -295 -1139
rect -353 -1207 -295 -1173
rect -353 -1241 -341 -1207
rect -307 -1241 -295 -1207
rect -353 -1275 -295 -1241
rect -353 -1309 -341 -1275
rect -307 -1309 -295 -1275
rect -353 -1343 -295 -1309
rect -353 -1377 -341 -1343
rect -307 -1377 -295 -1343
rect -353 -1411 -295 -1377
rect -353 -1445 -341 -1411
rect -307 -1445 -295 -1411
rect -353 -1479 -295 -1445
rect -353 -1513 -341 -1479
rect -307 -1513 -295 -1479
rect -353 -1547 -295 -1513
rect -353 -1581 -341 -1547
rect -307 -1581 -295 -1547
rect -353 -1615 -295 -1581
rect -353 -1649 -341 -1615
rect -307 -1649 -295 -1615
rect -353 -1683 -295 -1649
rect -353 -1717 -341 -1683
rect -307 -1717 -295 -1683
rect -353 -1751 -295 -1717
rect -353 -1785 -341 -1751
rect -307 -1785 -295 -1751
rect -353 -1819 -295 -1785
rect -353 -1853 -341 -1819
rect -307 -1853 -295 -1819
rect -353 -1887 -295 -1853
rect -353 -1921 -341 -1887
rect -307 -1921 -295 -1887
rect -353 -1955 -295 -1921
rect -353 -1989 -341 -1955
rect -307 -1989 -295 -1955
rect -353 -2023 -295 -1989
rect -353 -2057 -341 -2023
rect -307 -2057 -295 -2023
rect -353 -2091 -295 -2057
rect -353 -2125 -341 -2091
rect -307 -2125 -295 -2091
rect -353 -2159 -295 -2125
rect -353 -2193 -341 -2159
rect -307 -2193 -295 -2159
rect -353 -2227 -295 -2193
rect -353 -2261 -341 -2227
rect -307 -2261 -295 -2227
rect -353 -2295 -295 -2261
rect -353 -2329 -341 -2295
rect -307 -2329 -295 -2295
rect -353 -2363 -295 -2329
rect -353 -2397 -341 -2363
rect -307 -2397 -295 -2363
rect -353 -2431 -295 -2397
rect -353 -2465 -341 -2431
rect -307 -2465 -295 -2431
rect -353 -2500 -295 -2465
rect -245 2465 -187 2500
rect -245 2431 -233 2465
rect -199 2431 -187 2465
rect -245 2397 -187 2431
rect -245 2363 -233 2397
rect -199 2363 -187 2397
rect -245 2329 -187 2363
rect -245 2295 -233 2329
rect -199 2295 -187 2329
rect -245 2261 -187 2295
rect -245 2227 -233 2261
rect -199 2227 -187 2261
rect -245 2193 -187 2227
rect -245 2159 -233 2193
rect -199 2159 -187 2193
rect -245 2125 -187 2159
rect -245 2091 -233 2125
rect -199 2091 -187 2125
rect -245 2057 -187 2091
rect -245 2023 -233 2057
rect -199 2023 -187 2057
rect -245 1989 -187 2023
rect -245 1955 -233 1989
rect -199 1955 -187 1989
rect -245 1921 -187 1955
rect -245 1887 -233 1921
rect -199 1887 -187 1921
rect -245 1853 -187 1887
rect -245 1819 -233 1853
rect -199 1819 -187 1853
rect -245 1785 -187 1819
rect -245 1751 -233 1785
rect -199 1751 -187 1785
rect -245 1717 -187 1751
rect -245 1683 -233 1717
rect -199 1683 -187 1717
rect -245 1649 -187 1683
rect -245 1615 -233 1649
rect -199 1615 -187 1649
rect -245 1581 -187 1615
rect -245 1547 -233 1581
rect -199 1547 -187 1581
rect -245 1513 -187 1547
rect -245 1479 -233 1513
rect -199 1479 -187 1513
rect -245 1445 -187 1479
rect -245 1411 -233 1445
rect -199 1411 -187 1445
rect -245 1377 -187 1411
rect -245 1343 -233 1377
rect -199 1343 -187 1377
rect -245 1309 -187 1343
rect -245 1275 -233 1309
rect -199 1275 -187 1309
rect -245 1241 -187 1275
rect -245 1207 -233 1241
rect -199 1207 -187 1241
rect -245 1173 -187 1207
rect -245 1139 -233 1173
rect -199 1139 -187 1173
rect -245 1105 -187 1139
rect -245 1071 -233 1105
rect -199 1071 -187 1105
rect -245 1037 -187 1071
rect -245 1003 -233 1037
rect -199 1003 -187 1037
rect -245 969 -187 1003
rect -245 935 -233 969
rect -199 935 -187 969
rect -245 901 -187 935
rect -245 867 -233 901
rect -199 867 -187 901
rect -245 833 -187 867
rect -245 799 -233 833
rect -199 799 -187 833
rect -245 765 -187 799
rect -245 731 -233 765
rect -199 731 -187 765
rect -245 697 -187 731
rect -245 663 -233 697
rect -199 663 -187 697
rect -245 629 -187 663
rect -245 595 -233 629
rect -199 595 -187 629
rect -245 561 -187 595
rect -245 527 -233 561
rect -199 527 -187 561
rect -245 493 -187 527
rect -245 459 -233 493
rect -199 459 -187 493
rect -245 425 -187 459
rect -245 391 -233 425
rect -199 391 -187 425
rect -245 357 -187 391
rect -245 323 -233 357
rect -199 323 -187 357
rect -245 289 -187 323
rect -245 255 -233 289
rect -199 255 -187 289
rect -245 221 -187 255
rect -245 187 -233 221
rect -199 187 -187 221
rect -245 153 -187 187
rect -245 119 -233 153
rect -199 119 -187 153
rect -245 85 -187 119
rect -245 51 -233 85
rect -199 51 -187 85
rect -245 17 -187 51
rect -245 -17 -233 17
rect -199 -17 -187 17
rect -245 -51 -187 -17
rect -245 -85 -233 -51
rect -199 -85 -187 -51
rect -245 -119 -187 -85
rect -245 -153 -233 -119
rect -199 -153 -187 -119
rect -245 -187 -187 -153
rect -245 -221 -233 -187
rect -199 -221 -187 -187
rect -245 -255 -187 -221
rect -245 -289 -233 -255
rect -199 -289 -187 -255
rect -245 -323 -187 -289
rect -245 -357 -233 -323
rect -199 -357 -187 -323
rect -245 -391 -187 -357
rect -245 -425 -233 -391
rect -199 -425 -187 -391
rect -245 -459 -187 -425
rect -245 -493 -233 -459
rect -199 -493 -187 -459
rect -245 -527 -187 -493
rect -245 -561 -233 -527
rect -199 -561 -187 -527
rect -245 -595 -187 -561
rect -245 -629 -233 -595
rect -199 -629 -187 -595
rect -245 -663 -187 -629
rect -245 -697 -233 -663
rect -199 -697 -187 -663
rect -245 -731 -187 -697
rect -245 -765 -233 -731
rect -199 -765 -187 -731
rect -245 -799 -187 -765
rect -245 -833 -233 -799
rect -199 -833 -187 -799
rect -245 -867 -187 -833
rect -245 -901 -233 -867
rect -199 -901 -187 -867
rect -245 -935 -187 -901
rect -245 -969 -233 -935
rect -199 -969 -187 -935
rect -245 -1003 -187 -969
rect -245 -1037 -233 -1003
rect -199 -1037 -187 -1003
rect -245 -1071 -187 -1037
rect -245 -1105 -233 -1071
rect -199 -1105 -187 -1071
rect -245 -1139 -187 -1105
rect -245 -1173 -233 -1139
rect -199 -1173 -187 -1139
rect -245 -1207 -187 -1173
rect -245 -1241 -233 -1207
rect -199 -1241 -187 -1207
rect -245 -1275 -187 -1241
rect -245 -1309 -233 -1275
rect -199 -1309 -187 -1275
rect -245 -1343 -187 -1309
rect -245 -1377 -233 -1343
rect -199 -1377 -187 -1343
rect -245 -1411 -187 -1377
rect -245 -1445 -233 -1411
rect -199 -1445 -187 -1411
rect -245 -1479 -187 -1445
rect -245 -1513 -233 -1479
rect -199 -1513 -187 -1479
rect -245 -1547 -187 -1513
rect -245 -1581 -233 -1547
rect -199 -1581 -187 -1547
rect -245 -1615 -187 -1581
rect -245 -1649 -233 -1615
rect -199 -1649 -187 -1615
rect -245 -1683 -187 -1649
rect -245 -1717 -233 -1683
rect -199 -1717 -187 -1683
rect -245 -1751 -187 -1717
rect -245 -1785 -233 -1751
rect -199 -1785 -187 -1751
rect -245 -1819 -187 -1785
rect -245 -1853 -233 -1819
rect -199 -1853 -187 -1819
rect -245 -1887 -187 -1853
rect -245 -1921 -233 -1887
rect -199 -1921 -187 -1887
rect -245 -1955 -187 -1921
rect -245 -1989 -233 -1955
rect -199 -1989 -187 -1955
rect -245 -2023 -187 -1989
rect -245 -2057 -233 -2023
rect -199 -2057 -187 -2023
rect -245 -2091 -187 -2057
rect -245 -2125 -233 -2091
rect -199 -2125 -187 -2091
rect -245 -2159 -187 -2125
rect -245 -2193 -233 -2159
rect -199 -2193 -187 -2159
rect -245 -2227 -187 -2193
rect -245 -2261 -233 -2227
rect -199 -2261 -187 -2227
rect -245 -2295 -187 -2261
rect -245 -2329 -233 -2295
rect -199 -2329 -187 -2295
rect -245 -2363 -187 -2329
rect -245 -2397 -233 -2363
rect -199 -2397 -187 -2363
rect -245 -2431 -187 -2397
rect -245 -2465 -233 -2431
rect -199 -2465 -187 -2431
rect -245 -2500 -187 -2465
rect -137 2465 -79 2500
rect -137 2431 -125 2465
rect -91 2431 -79 2465
rect -137 2397 -79 2431
rect -137 2363 -125 2397
rect -91 2363 -79 2397
rect -137 2329 -79 2363
rect -137 2295 -125 2329
rect -91 2295 -79 2329
rect -137 2261 -79 2295
rect -137 2227 -125 2261
rect -91 2227 -79 2261
rect -137 2193 -79 2227
rect -137 2159 -125 2193
rect -91 2159 -79 2193
rect -137 2125 -79 2159
rect -137 2091 -125 2125
rect -91 2091 -79 2125
rect -137 2057 -79 2091
rect -137 2023 -125 2057
rect -91 2023 -79 2057
rect -137 1989 -79 2023
rect -137 1955 -125 1989
rect -91 1955 -79 1989
rect -137 1921 -79 1955
rect -137 1887 -125 1921
rect -91 1887 -79 1921
rect -137 1853 -79 1887
rect -137 1819 -125 1853
rect -91 1819 -79 1853
rect -137 1785 -79 1819
rect -137 1751 -125 1785
rect -91 1751 -79 1785
rect -137 1717 -79 1751
rect -137 1683 -125 1717
rect -91 1683 -79 1717
rect -137 1649 -79 1683
rect -137 1615 -125 1649
rect -91 1615 -79 1649
rect -137 1581 -79 1615
rect -137 1547 -125 1581
rect -91 1547 -79 1581
rect -137 1513 -79 1547
rect -137 1479 -125 1513
rect -91 1479 -79 1513
rect -137 1445 -79 1479
rect -137 1411 -125 1445
rect -91 1411 -79 1445
rect -137 1377 -79 1411
rect -137 1343 -125 1377
rect -91 1343 -79 1377
rect -137 1309 -79 1343
rect -137 1275 -125 1309
rect -91 1275 -79 1309
rect -137 1241 -79 1275
rect -137 1207 -125 1241
rect -91 1207 -79 1241
rect -137 1173 -79 1207
rect -137 1139 -125 1173
rect -91 1139 -79 1173
rect -137 1105 -79 1139
rect -137 1071 -125 1105
rect -91 1071 -79 1105
rect -137 1037 -79 1071
rect -137 1003 -125 1037
rect -91 1003 -79 1037
rect -137 969 -79 1003
rect -137 935 -125 969
rect -91 935 -79 969
rect -137 901 -79 935
rect -137 867 -125 901
rect -91 867 -79 901
rect -137 833 -79 867
rect -137 799 -125 833
rect -91 799 -79 833
rect -137 765 -79 799
rect -137 731 -125 765
rect -91 731 -79 765
rect -137 697 -79 731
rect -137 663 -125 697
rect -91 663 -79 697
rect -137 629 -79 663
rect -137 595 -125 629
rect -91 595 -79 629
rect -137 561 -79 595
rect -137 527 -125 561
rect -91 527 -79 561
rect -137 493 -79 527
rect -137 459 -125 493
rect -91 459 -79 493
rect -137 425 -79 459
rect -137 391 -125 425
rect -91 391 -79 425
rect -137 357 -79 391
rect -137 323 -125 357
rect -91 323 -79 357
rect -137 289 -79 323
rect -137 255 -125 289
rect -91 255 -79 289
rect -137 221 -79 255
rect -137 187 -125 221
rect -91 187 -79 221
rect -137 153 -79 187
rect -137 119 -125 153
rect -91 119 -79 153
rect -137 85 -79 119
rect -137 51 -125 85
rect -91 51 -79 85
rect -137 17 -79 51
rect -137 -17 -125 17
rect -91 -17 -79 17
rect -137 -51 -79 -17
rect -137 -85 -125 -51
rect -91 -85 -79 -51
rect -137 -119 -79 -85
rect -137 -153 -125 -119
rect -91 -153 -79 -119
rect -137 -187 -79 -153
rect -137 -221 -125 -187
rect -91 -221 -79 -187
rect -137 -255 -79 -221
rect -137 -289 -125 -255
rect -91 -289 -79 -255
rect -137 -323 -79 -289
rect -137 -357 -125 -323
rect -91 -357 -79 -323
rect -137 -391 -79 -357
rect -137 -425 -125 -391
rect -91 -425 -79 -391
rect -137 -459 -79 -425
rect -137 -493 -125 -459
rect -91 -493 -79 -459
rect -137 -527 -79 -493
rect -137 -561 -125 -527
rect -91 -561 -79 -527
rect -137 -595 -79 -561
rect -137 -629 -125 -595
rect -91 -629 -79 -595
rect -137 -663 -79 -629
rect -137 -697 -125 -663
rect -91 -697 -79 -663
rect -137 -731 -79 -697
rect -137 -765 -125 -731
rect -91 -765 -79 -731
rect -137 -799 -79 -765
rect -137 -833 -125 -799
rect -91 -833 -79 -799
rect -137 -867 -79 -833
rect -137 -901 -125 -867
rect -91 -901 -79 -867
rect -137 -935 -79 -901
rect -137 -969 -125 -935
rect -91 -969 -79 -935
rect -137 -1003 -79 -969
rect -137 -1037 -125 -1003
rect -91 -1037 -79 -1003
rect -137 -1071 -79 -1037
rect -137 -1105 -125 -1071
rect -91 -1105 -79 -1071
rect -137 -1139 -79 -1105
rect -137 -1173 -125 -1139
rect -91 -1173 -79 -1139
rect -137 -1207 -79 -1173
rect -137 -1241 -125 -1207
rect -91 -1241 -79 -1207
rect -137 -1275 -79 -1241
rect -137 -1309 -125 -1275
rect -91 -1309 -79 -1275
rect -137 -1343 -79 -1309
rect -137 -1377 -125 -1343
rect -91 -1377 -79 -1343
rect -137 -1411 -79 -1377
rect -137 -1445 -125 -1411
rect -91 -1445 -79 -1411
rect -137 -1479 -79 -1445
rect -137 -1513 -125 -1479
rect -91 -1513 -79 -1479
rect -137 -1547 -79 -1513
rect -137 -1581 -125 -1547
rect -91 -1581 -79 -1547
rect -137 -1615 -79 -1581
rect -137 -1649 -125 -1615
rect -91 -1649 -79 -1615
rect -137 -1683 -79 -1649
rect -137 -1717 -125 -1683
rect -91 -1717 -79 -1683
rect -137 -1751 -79 -1717
rect -137 -1785 -125 -1751
rect -91 -1785 -79 -1751
rect -137 -1819 -79 -1785
rect -137 -1853 -125 -1819
rect -91 -1853 -79 -1819
rect -137 -1887 -79 -1853
rect -137 -1921 -125 -1887
rect -91 -1921 -79 -1887
rect -137 -1955 -79 -1921
rect -137 -1989 -125 -1955
rect -91 -1989 -79 -1955
rect -137 -2023 -79 -1989
rect -137 -2057 -125 -2023
rect -91 -2057 -79 -2023
rect -137 -2091 -79 -2057
rect -137 -2125 -125 -2091
rect -91 -2125 -79 -2091
rect -137 -2159 -79 -2125
rect -137 -2193 -125 -2159
rect -91 -2193 -79 -2159
rect -137 -2227 -79 -2193
rect -137 -2261 -125 -2227
rect -91 -2261 -79 -2227
rect -137 -2295 -79 -2261
rect -137 -2329 -125 -2295
rect -91 -2329 -79 -2295
rect -137 -2363 -79 -2329
rect -137 -2397 -125 -2363
rect -91 -2397 -79 -2363
rect -137 -2431 -79 -2397
rect -137 -2465 -125 -2431
rect -91 -2465 -79 -2431
rect -137 -2500 -79 -2465
rect -29 2465 29 2500
rect -29 2431 -17 2465
rect 17 2431 29 2465
rect -29 2397 29 2431
rect -29 2363 -17 2397
rect 17 2363 29 2397
rect -29 2329 29 2363
rect -29 2295 -17 2329
rect 17 2295 29 2329
rect -29 2261 29 2295
rect -29 2227 -17 2261
rect 17 2227 29 2261
rect -29 2193 29 2227
rect -29 2159 -17 2193
rect 17 2159 29 2193
rect -29 2125 29 2159
rect -29 2091 -17 2125
rect 17 2091 29 2125
rect -29 2057 29 2091
rect -29 2023 -17 2057
rect 17 2023 29 2057
rect -29 1989 29 2023
rect -29 1955 -17 1989
rect 17 1955 29 1989
rect -29 1921 29 1955
rect -29 1887 -17 1921
rect 17 1887 29 1921
rect -29 1853 29 1887
rect -29 1819 -17 1853
rect 17 1819 29 1853
rect -29 1785 29 1819
rect -29 1751 -17 1785
rect 17 1751 29 1785
rect -29 1717 29 1751
rect -29 1683 -17 1717
rect 17 1683 29 1717
rect -29 1649 29 1683
rect -29 1615 -17 1649
rect 17 1615 29 1649
rect -29 1581 29 1615
rect -29 1547 -17 1581
rect 17 1547 29 1581
rect -29 1513 29 1547
rect -29 1479 -17 1513
rect 17 1479 29 1513
rect -29 1445 29 1479
rect -29 1411 -17 1445
rect 17 1411 29 1445
rect -29 1377 29 1411
rect -29 1343 -17 1377
rect 17 1343 29 1377
rect -29 1309 29 1343
rect -29 1275 -17 1309
rect 17 1275 29 1309
rect -29 1241 29 1275
rect -29 1207 -17 1241
rect 17 1207 29 1241
rect -29 1173 29 1207
rect -29 1139 -17 1173
rect 17 1139 29 1173
rect -29 1105 29 1139
rect -29 1071 -17 1105
rect 17 1071 29 1105
rect -29 1037 29 1071
rect -29 1003 -17 1037
rect 17 1003 29 1037
rect -29 969 29 1003
rect -29 935 -17 969
rect 17 935 29 969
rect -29 901 29 935
rect -29 867 -17 901
rect 17 867 29 901
rect -29 833 29 867
rect -29 799 -17 833
rect 17 799 29 833
rect -29 765 29 799
rect -29 731 -17 765
rect 17 731 29 765
rect -29 697 29 731
rect -29 663 -17 697
rect 17 663 29 697
rect -29 629 29 663
rect -29 595 -17 629
rect 17 595 29 629
rect -29 561 29 595
rect -29 527 -17 561
rect 17 527 29 561
rect -29 493 29 527
rect -29 459 -17 493
rect 17 459 29 493
rect -29 425 29 459
rect -29 391 -17 425
rect 17 391 29 425
rect -29 357 29 391
rect -29 323 -17 357
rect 17 323 29 357
rect -29 289 29 323
rect -29 255 -17 289
rect 17 255 29 289
rect -29 221 29 255
rect -29 187 -17 221
rect 17 187 29 221
rect -29 153 29 187
rect -29 119 -17 153
rect 17 119 29 153
rect -29 85 29 119
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -119 29 -85
rect -29 -153 -17 -119
rect 17 -153 29 -119
rect -29 -187 29 -153
rect -29 -221 -17 -187
rect 17 -221 29 -187
rect -29 -255 29 -221
rect -29 -289 -17 -255
rect 17 -289 29 -255
rect -29 -323 29 -289
rect -29 -357 -17 -323
rect 17 -357 29 -323
rect -29 -391 29 -357
rect -29 -425 -17 -391
rect 17 -425 29 -391
rect -29 -459 29 -425
rect -29 -493 -17 -459
rect 17 -493 29 -459
rect -29 -527 29 -493
rect -29 -561 -17 -527
rect 17 -561 29 -527
rect -29 -595 29 -561
rect -29 -629 -17 -595
rect 17 -629 29 -595
rect -29 -663 29 -629
rect -29 -697 -17 -663
rect 17 -697 29 -663
rect -29 -731 29 -697
rect -29 -765 -17 -731
rect 17 -765 29 -731
rect -29 -799 29 -765
rect -29 -833 -17 -799
rect 17 -833 29 -799
rect -29 -867 29 -833
rect -29 -901 -17 -867
rect 17 -901 29 -867
rect -29 -935 29 -901
rect -29 -969 -17 -935
rect 17 -969 29 -935
rect -29 -1003 29 -969
rect -29 -1037 -17 -1003
rect 17 -1037 29 -1003
rect -29 -1071 29 -1037
rect -29 -1105 -17 -1071
rect 17 -1105 29 -1071
rect -29 -1139 29 -1105
rect -29 -1173 -17 -1139
rect 17 -1173 29 -1139
rect -29 -1207 29 -1173
rect -29 -1241 -17 -1207
rect 17 -1241 29 -1207
rect -29 -1275 29 -1241
rect -29 -1309 -17 -1275
rect 17 -1309 29 -1275
rect -29 -1343 29 -1309
rect -29 -1377 -17 -1343
rect 17 -1377 29 -1343
rect -29 -1411 29 -1377
rect -29 -1445 -17 -1411
rect 17 -1445 29 -1411
rect -29 -1479 29 -1445
rect -29 -1513 -17 -1479
rect 17 -1513 29 -1479
rect -29 -1547 29 -1513
rect -29 -1581 -17 -1547
rect 17 -1581 29 -1547
rect -29 -1615 29 -1581
rect -29 -1649 -17 -1615
rect 17 -1649 29 -1615
rect -29 -1683 29 -1649
rect -29 -1717 -17 -1683
rect 17 -1717 29 -1683
rect -29 -1751 29 -1717
rect -29 -1785 -17 -1751
rect 17 -1785 29 -1751
rect -29 -1819 29 -1785
rect -29 -1853 -17 -1819
rect 17 -1853 29 -1819
rect -29 -1887 29 -1853
rect -29 -1921 -17 -1887
rect 17 -1921 29 -1887
rect -29 -1955 29 -1921
rect -29 -1989 -17 -1955
rect 17 -1989 29 -1955
rect -29 -2023 29 -1989
rect -29 -2057 -17 -2023
rect 17 -2057 29 -2023
rect -29 -2091 29 -2057
rect -29 -2125 -17 -2091
rect 17 -2125 29 -2091
rect -29 -2159 29 -2125
rect -29 -2193 -17 -2159
rect 17 -2193 29 -2159
rect -29 -2227 29 -2193
rect -29 -2261 -17 -2227
rect 17 -2261 29 -2227
rect -29 -2295 29 -2261
rect -29 -2329 -17 -2295
rect 17 -2329 29 -2295
rect -29 -2363 29 -2329
rect -29 -2397 -17 -2363
rect 17 -2397 29 -2363
rect -29 -2431 29 -2397
rect -29 -2465 -17 -2431
rect 17 -2465 29 -2431
rect -29 -2500 29 -2465
rect 79 2465 137 2500
rect 79 2431 91 2465
rect 125 2431 137 2465
rect 79 2397 137 2431
rect 79 2363 91 2397
rect 125 2363 137 2397
rect 79 2329 137 2363
rect 79 2295 91 2329
rect 125 2295 137 2329
rect 79 2261 137 2295
rect 79 2227 91 2261
rect 125 2227 137 2261
rect 79 2193 137 2227
rect 79 2159 91 2193
rect 125 2159 137 2193
rect 79 2125 137 2159
rect 79 2091 91 2125
rect 125 2091 137 2125
rect 79 2057 137 2091
rect 79 2023 91 2057
rect 125 2023 137 2057
rect 79 1989 137 2023
rect 79 1955 91 1989
rect 125 1955 137 1989
rect 79 1921 137 1955
rect 79 1887 91 1921
rect 125 1887 137 1921
rect 79 1853 137 1887
rect 79 1819 91 1853
rect 125 1819 137 1853
rect 79 1785 137 1819
rect 79 1751 91 1785
rect 125 1751 137 1785
rect 79 1717 137 1751
rect 79 1683 91 1717
rect 125 1683 137 1717
rect 79 1649 137 1683
rect 79 1615 91 1649
rect 125 1615 137 1649
rect 79 1581 137 1615
rect 79 1547 91 1581
rect 125 1547 137 1581
rect 79 1513 137 1547
rect 79 1479 91 1513
rect 125 1479 137 1513
rect 79 1445 137 1479
rect 79 1411 91 1445
rect 125 1411 137 1445
rect 79 1377 137 1411
rect 79 1343 91 1377
rect 125 1343 137 1377
rect 79 1309 137 1343
rect 79 1275 91 1309
rect 125 1275 137 1309
rect 79 1241 137 1275
rect 79 1207 91 1241
rect 125 1207 137 1241
rect 79 1173 137 1207
rect 79 1139 91 1173
rect 125 1139 137 1173
rect 79 1105 137 1139
rect 79 1071 91 1105
rect 125 1071 137 1105
rect 79 1037 137 1071
rect 79 1003 91 1037
rect 125 1003 137 1037
rect 79 969 137 1003
rect 79 935 91 969
rect 125 935 137 969
rect 79 901 137 935
rect 79 867 91 901
rect 125 867 137 901
rect 79 833 137 867
rect 79 799 91 833
rect 125 799 137 833
rect 79 765 137 799
rect 79 731 91 765
rect 125 731 137 765
rect 79 697 137 731
rect 79 663 91 697
rect 125 663 137 697
rect 79 629 137 663
rect 79 595 91 629
rect 125 595 137 629
rect 79 561 137 595
rect 79 527 91 561
rect 125 527 137 561
rect 79 493 137 527
rect 79 459 91 493
rect 125 459 137 493
rect 79 425 137 459
rect 79 391 91 425
rect 125 391 137 425
rect 79 357 137 391
rect 79 323 91 357
rect 125 323 137 357
rect 79 289 137 323
rect 79 255 91 289
rect 125 255 137 289
rect 79 221 137 255
rect 79 187 91 221
rect 125 187 137 221
rect 79 153 137 187
rect 79 119 91 153
rect 125 119 137 153
rect 79 85 137 119
rect 79 51 91 85
rect 125 51 137 85
rect 79 17 137 51
rect 79 -17 91 17
rect 125 -17 137 17
rect 79 -51 137 -17
rect 79 -85 91 -51
rect 125 -85 137 -51
rect 79 -119 137 -85
rect 79 -153 91 -119
rect 125 -153 137 -119
rect 79 -187 137 -153
rect 79 -221 91 -187
rect 125 -221 137 -187
rect 79 -255 137 -221
rect 79 -289 91 -255
rect 125 -289 137 -255
rect 79 -323 137 -289
rect 79 -357 91 -323
rect 125 -357 137 -323
rect 79 -391 137 -357
rect 79 -425 91 -391
rect 125 -425 137 -391
rect 79 -459 137 -425
rect 79 -493 91 -459
rect 125 -493 137 -459
rect 79 -527 137 -493
rect 79 -561 91 -527
rect 125 -561 137 -527
rect 79 -595 137 -561
rect 79 -629 91 -595
rect 125 -629 137 -595
rect 79 -663 137 -629
rect 79 -697 91 -663
rect 125 -697 137 -663
rect 79 -731 137 -697
rect 79 -765 91 -731
rect 125 -765 137 -731
rect 79 -799 137 -765
rect 79 -833 91 -799
rect 125 -833 137 -799
rect 79 -867 137 -833
rect 79 -901 91 -867
rect 125 -901 137 -867
rect 79 -935 137 -901
rect 79 -969 91 -935
rect 125 -969 137 -935
rect 79 -1003 137 -969
rect 79 -1037 91 -1003
rect 125 -1037 137 -1003
rect 79 -1071 137 -1037
rect 79 -1105 91 -1071
rect 125 -1105 137 -1071
rect 79 -1139 137 -1105
rect 79 -1173 91 -1139
rect 125 -1173 137 -1139
rect 79 -1207 137 -1173
rect 79 -1241 91 -1207
rect 125 -1241 137 -1207
rect 79 -1275 137 -1241
rect 79 -1309 91 -1275
rect 125 -1309 137 -1275
rect 79 -1343 137 -1309
rect 79 -1377 91 -1343
rect 125 -1377 137 -1343
rect 79 -1411 137 -1377
rect 79 -1445 91 -1411
rect 125 -1445 137 -1411
rect 79 -1479 137 -1445
rect 79 -1513 91 -1479
rect 125 -1513 137 -1479
rect 79 -1547 137 -1513
rect 79 -1581 91 -1547
rect 125 -1581 137 -1547
rect 79 -1615 137 -1581
rect 79 -1649 91 -1615
rect 125 -1649 137 -1615
rect 79 -1683 137 -1649
rect 79 -1717 91 -1683
rect 125 -1717 137 -1683
rect 79 -1751 137 -1717
rect 79 -1785 91 -1751
rect 125 -1785 137 -1751
rect 79 -1819 137 -1785
rect 79 -1853 91 -1819
rect 125 -1853 137 -1819
rect 79 -1887 137 -1853
rect 79 -1921 91 -1887
rect 125 -1921 137 -1887
rect 79 -1955 137 -1921
rect 79 -1989 91 -1955
rect 125 -1989 137 -1955
rect 79 -2023 137 -1989
rect 79 -2057 91 -2023
rect 125 -2057 137 -2023
rect 79 -2091 137 -2057
rect 79 -2125 91 -2091
rect 125 -2125 137 -2091
rect 79 -2159 137 -2125
rect 79 -2193 91 -2159
rect 125 -2193 137 -2159
rect 79 -2227 137 -2193
rect 79 -2261 91 -2227
rect 125 -2261 137 -2227
rect 79 -2295 137 -2261
rect 79 -2329 91 -2295
rect 125 -2329 137 -2295
rect 79 -2363 137 -2329
rect 79 -2397 91 -2363
rect 125 -2397 137 -2363
rect 79 -2431 137 -2397
rect 79 -2465 91 -2431
rect 125 -2465 137 -2431
rect 79 -2500 137 -2465
rect 187 2465 245 2500
rect 187 2431 199 2465
rect 233 2431 245 2465
rect 187 2397 245 2431
rect 187 2363 199 2397
rect 233 2363 245 2397
rect 187 2329 245 2363
rect 187 2295 199 2329
rect 233 2295 245 2329
rect 187 2261 245 2295
rect 187 2227 199 2261
rect 233 2227 245 2261
rect 187 2193 245 2227
rect 187 2159 199 2193
rect 233 2159 245 2193
rect 187 2125 245 2159
rect 187 2091 199 2125
rect 233 2091 245 2125
rect 187 2057 245 2091
rect 187 2023 199 2057
rect 233 2023 245 2057
rect 187 1989 245 2023
rect 187 1955 199 1989
rect 233 1955 245 1989
rect 187 1921 245 1955
rect 187 1887 199 1921
rect 233 1887 245 1921
rect 187 1853 245 1887
rect 187 1819 199 1853
rect 233 1819 245 1853
rect 187 1785 245 1819
rect 187 1751 199 1785
rect 233 1751 245 1785
rect 187 1717 245 1751
rect 187 1683 199 1717
rect 233 1683 245 1717
rect 187 1649 245 1683
rect 187 1615 199 1649
rect 233 1615 245 1649
rect 187 1581 245 1615
rect 187 1547 199 1581
rect 233 1547 245 1581
rect 187 1513 245 1547
rect 187 1479 199 1513
rect 233 1479 245 1513
rect 187 1445 245 1479
rect 187 1411 199 1445
rect 233 1411 245 1445
rect 187 1377 245 1411
rect 187 1343 199 1377
rect 233 1343 245 1377
rect 187 1309 245 1343
rect 187 1275 199 1309
rect 233 1275 245 1309
rect 187 1241 245 1275
rect 187 1207 199 1241
rect 233 1207 245 1241
rect 187 1173 245 1207
rect 187 1139 199 1173
rect 233 1139 245 1173
rect 187 1105 245 1139
rect 187 1071 199 1105
rect 233 1071 245 1105
rect 187 1037 245 1071
rect 187 1003 199 1037
rect 233 1003 245 1037
rect 187 969 245 1003
rect 187 935 199 969
rect 233 935 245 969
rect 187 901 245 935
rect 187 867 199 901
rect 233 867 245 901
rect 187 833 245 867
rect 187 799 199 833
rect 233 799 245 833
rect 187 765 245 799
rect 187 731 199 765
rect 233 731 245 765
rect 187 697 245 731
rect 187 663 199 697
rect 233 663 245 697
rect 187 629 245 663
rect 187 595 199 629
rect 233 595 245 629
rect 187 561 245 595
rect 187 527 199 561
rect 233 527 245 561
rect 187 493 245 527
rect 187 459 199 493
rect 233 459 245 493
rect 187 425 245 459
rect 187 391 199 425
rect 233 391 245 425
rect 187 357 245 391
rect 187 323 199 357
rect 233 323 245 357
rect 187 289 245 323
rect 187 255 199 289
rect 233 255 245 289
rect 187 221 245 255
rect 187 187 199 221
rect 233 187 245 221
rect 187 153 245 187
rect 187 119 199 153
rect 233 119 245 153
rect 187 85 245 119
rect 187 51 199 85
rect 233 51 245 85
rect 187 17 245 51
rect 187 -17 199 17
rect 233 -17 245 17
rect 187 -51 245 -17
rect 187 -85 199 -51
rect 233 -85 245 -51
rect 187 -119 245 -85
rect 187 -153 199 -119
rect 233 -153 245 -119
rect 187 -187 245 -153
rect 187 -221 199 -187
rect 233 -221 245 -187
rect 187 -255 245 -221
rect 187 -289 199 -255
rect 233 -289 245 -255
rect 187 -323 245 -289
rect 187 -357 199 -323
rect 233 -357 245 -323
rect 187 -391 245 -357
rect 187 -425 199 -391
rect 233 -425 245 -391
rect 187 -459 245 -425
rect 187 -493 199 -459
rect 233 -493 245 -459
rect 187 -527 245 -493
rect 187 -561 199 -527
rect 233 -561 245 -527
rect 187 -595 245 -561
rect 187 -629 199 -595
rect 233 -629 245 -595
rect 187 -663 245 -629
rect 187 -697 199 -663
rect 233 -697 245 -663
rect 187 -731 245 -697
rect 187 -765 199 -731
rect 233 -765 245 -731
rect 187 -799 245 -765
rect 187 -833 199 -799
rect 233 -833 245 -799
rect 187 -867 245 -833
rect 187 -901 199 -867
rect 233 -901 245 -867
rect 187 -935 245 -901
rect 187 -969 199 -935
rect 233 -969 245 -935
rect 187 -1003 245 -969
rect 187 -1037 199 -1003
rect 233 -1037 245 -1003
rect 187 -1071 245 -1037
rect 187 -1105 199 -1071
rect 233 -1105 245 -1071
rect 187 -1139 245 -1105
rect 187 -1173 199 -1139
rect 233 -1173 245 -1139
rect 187 -1207 245 -1173
rect 187 -1241 199 -1207
rect 233 -1241 245 -1207
rect 187 -1275 245 -1241
rect 187 -1309 199 -1275
rect 233 -1309 245 -1275
rect 187 -1343 245 -1309
rect 187 -1377 199 -1343
rect 233 -1377 245 -1343
rect 187 -1411 245 -1377
rect 187 -1445 199 -1411
rect 233 -1445 245 -1411
rect 187 -1479 245 -1445
rect 187 -1513 199 -1479
rect 233 -1513 245 -1479
rect 187 -1547 245 -1513
rect 187 -1581 199 -1547
rect 233 -1581 245 -1547
rect 187 -1615 245 -1581
rect 187 -1649 199 -1615
rect 233 -1649 245 -1615
rect 187 -1683 245 -1649
rect 187 -1717 199 -1683
rect 233 -1717 245 -1683
rect 187 -1751 245 -1717
rect 187 -1785 199 -1751
rect 233 -1785 245 -1751
rect 187 -1819 245 -1785
rect 187 -1853 199 -1819
rect 233 -1853 245 -1819
rect 187 -1887 245 -1853
rect 187 -1921 199 -1887
rect 233 -1921 245 -1887
rect 187 -1955 245 -1921
rect 187 -1989 199 -1955
rect 233 -1989 245 -1955
rect 187 -2023 245 -1989
rect 187 -2057 199 -2023
rect 233 -2057 245 -2023
rect 187 -2091 245 -2057
rect 187 -2125 199 -2091
rect 233 -2125 245 -2091
rect 187 -2159 245 -2125
rect 187 -2193 199 -2159
rect 233 -2193 245 -2159
rect 187 -2227 245 -2193
rect 187 -2261 199 -2227
rect 233 -2261 245 -2227
rect 187 -2295 245 -2261
rect 187 -2329 199 -2295
rect 233 -2329 245 -2295
rect 187 -2363 245 -2329
rect 187 -2397 199 -2363
rect 233 -2397 245 -2363
rect 187 -2431 245 -2397
rect 187 -2465 199 -2431
rect 233 -2465 245 -2431
rect 187 -2500 245 -2465
rect 295 2465 353 2500
rect 295 2431 307 2465
rect 341 2431 353 2465
rect 295 2397 353 2431
rect 295 2363 307 2397
rect 341 2363 353 2397
rect 295 2329 353 2363
rect 295 2295 307 2329
rect 341 2295 353 2329
rect 295 2261 353 2295
rect 295 2227 307 2261
rect 341 2227 353 2261
rect 295 2193 353 2227
rect 295 2159 307 2193
rect 341 2159 353 2193
rect 295 2125 353 2159
rect 295 2091 307 2125
rect 341 2091 353 2125
rect 295 2057 353 2091
rect 295 2023 307 2057
rect 341 2023 353 2057
rect 295 1989 353 2023
rect 295 1955 307 1989
rect 341 1955 353 1989
rect 295 1921 353 1955
rect 295 1887 307 1921
rect 341 1887 353 1921
rect 295 1853 353 1887
rect 295 1819 307 1853
rect 341 1819 353 1853
rect 295 1785 353 1819
rect 295 1751 307 1785
rect 341 1751 353 1785
rect 295 1717 353 1751
rect 295 1683 307 1717
rect 341 1683 353 1717
rect 295 1649 353 1683
rect 295 1615 307 1649
rect 341 1615 353 1649
rect 295 1581 353 1615
rect 295 1547 307 1581
rect 341 1547 353 1581
rect 295 1513 353 1547
rect 295 1479 307 1513
rect 341 1479 353 1513
rect 295 1445 353 1479
rect 295 1411 307 1445
rect 341 1411 353 1445
rect 295 1377 353 1411
rect 295 1343 307 1377
rect 341 1343 353 1377
rect 295 1309 353 1343
rect 295 1275 307 1309
rect 341 1275 353 1309
rect 295 1241 353 1275
rect 295 1207 307 1241
rect 341 1207 353 1241
rect 295 1173 353 1207
rect 295 1139 307 1173
rect 341 1139 353 1173
rect 295 1105 353 1139
rect 295 1071 307 1105
rect 341 1071 353 1105
rect 295 1037 353 1071
rect 295 1003 307 1037
rect 341 1003 353 1037
rect 295 969 353 1003
rect 295 935 307 969
rect 341 935 353 969
rect 295 901 353 935
rect 295 867 307 901
rect 341 867 353 901
rect 295 833 353 867
rect 295 799 307 833
rect 341 799 353 833
rect 295 765 353 799
rect 295 731 307 765
rect 341 731 353 765
rect 295 697 353 731
rect 295 663 307 697
rect 341 663 353 697
rect 295 629 353 663
rect 295 595 307 629
rect 341 595 353 629
rect 295 561 353 595
rect 295 527 307 561
rect 341 527 353 561
rect 295 493 353 527
rect 295 459 307 493
rect 341 459 353 493
rect 295 425 353 459
rect 295 391 307 425
rect 341 391 353 425
rect 295 357 353 391
rect 295 323 307 357
rect 341 323 353 357
rect 295 289 353 323
rect 295 255 307 289
rect 341 255 353 289
rect 295 221 353 255
rect 295 187 307 221
rect 341 187 353 221
rect 295 153 353 187
rect 295 119 307 153
rect 341 119 353 153
rect 295 85 353 119
rect 295 51 307 85
rect 341 51 353 85
rect 295 17 353 51
rect 295 -17 307 17
rect 341 -17 353 17
rect 295 -51 353 -17
rect 295 -85 307 -51
rect 341 -85 353 -51
rect 295 -119 353 -85
rect 295 -153 307 -119
rect 341 -153 353 -119
rect 295 -187 353 -153
rect 295 -221 307 -187
rect 341 -221 353 -187
rect 295 -255 353 -221
rect 295 -289 307 -255
rect 341 -289 353 -255
rect 295 -323 353 -289
rect 295 -357 307 -323
rect 341 -357 353 -323
rect 295 -391 353 -357
rect 295 -425 307 -391
rect 341 -425 353 -391
rect 295 -459 353 -425
rect 295 -493 307 -459
rect 341 -493 353 -459
rect 295 -527 353 -493
rect 295 -561 307 -527
rect 341 -561 353 -527
rect 295 -595 353 -561
rect 295 -629 307 -595
rect 341 -629 353 -595
rect 295 -663 353 -629
rect 295 -697 307 -663
rect 341 -697 353 -663
rect 295 -731 353 -697
rect 295 -765 307 -731
rect 341 -765 353 -731
rect 295 -799 353 -765
rect 295 -833 307 -799
rect 341 -833 353 -799
rect 295 -867 353 -833
rect 295 -901 307 -867
rect 341 -901 353 -867
rect 295 -935 353 -901
rect 295 -969 307 -935
rect 341 -969 353 -935
rect 295 -1003 353 -969
rect 295 -1037 307 -1003
rect 341 -1037 353 -1003
rect 295 -1071 353 -1037
rect 295 -1105 307 -1071
rect 341 -1105 353 -1071
rect 295 -1139 353 -1105
rect 295 -1173 307 -1139
rect 341 -1173 353 -1139
rect 295 -1207 353 -1173
rect 295 -1241 307 -1207
rect 341 -1241 353 -1207
rect 295 -1275 353 -1241
rect 295 -1309 307 -1275
rect 341 -1309 353 -1275
rect 295 -1343 353 -1309
rect 295 -1377 307 -1343
rect 341 -1377 353 -1343
rect 295 -1411 353 -1377
rect 295 -1445 307 -1411
rect 341 -1445 353 -1411
rect 295 -1479 353 -1445
rect 295 -1513 307 -1479
rect 341 -1513 353 -1479
rect 295 -1547 353 -1513
rect 295 -1581 307 -1547
rect 341 -1581 353 -1547
rect 295 -1615 353 -1581
rect 295 -1649 307 -1615
rect 341 -1649 353 -1615
rect 295 -1683 353 -1649
rect 295 -1717 307 -1683
rect 341 -1717 353 -1683
rect 295 -1751 353 -1717
rect 295 -1785 307 -1751
rect 341 -1785 353 -1751
rect 295 -1819 353 -1785
rect 295 -1853 307 -1819
rect 341 -1853 353 -1819
rect 295 -1887 353 -1853
rect 295 -1921 307 -1887
rect 341 -1921 353 -1887
rect 295 -1955 353 -1921
rect 295 -1989 307 -1955
rect 341 -1989 353 -1955
rect 295 -2023 353 -1989
rect 295 -2057 307 -2023
rect 341 -2057 353 -2023
rect 295 -2091 353 -2057
rect 295 -2125 307 -2091
rect 341 -2125 353 -2091
rect 295 -2159 353 -2125
rect 295 -2193 307 -2159
rect 341 -2193 353 -2159
rect 295 -2227 353 -2193
rect 295 -2261 307 -2227
rect 341 -2261 353 -2227
rect 295 -2295 353 -2261
rect 295 -2329 307 -2295
rect 341 -2329 353 -2295
rect 295 -2363 353 -2329
rect 295 -2397 307 -2363
rect 341 -2397 353 -2363
rect 295 -2431 353 -2397
rect 295 -2465 307 -2431
rect 341 -2465 353 -2431
rect 295 -2500 353 -2465
rect 403 2465 461 2500
rect 403 2431 415 2465
rect 449 2431 461 2465
rect 403 2397 461 2431
rect 403 2363 415 2397
rect 449 2363 461 2397
rect 403 2329 461 2363
rect 403 2295 415 2329
rect 449 2295 461 2329
rect 403 2261 461 2295
rect 403 2227 415 2261
rect 449 2227 461 2261
rect 403 2193 461 2227
rect 403 2159 415 2193
rect 449 2159 461 2193
rect 403 2125 461 2159
rect 403 2091 415 2125
rect 449 2091 461 2125
rect 403 2057 461 2091
rect 403 2023 415 2057
rect 449 2023 461 2057
rect 403 1989 461 2023
rect 403 1955 415 1989
rect 449 1955 461 1989
rect 403 1921 461 1955
rect 403 1887 415 1921
rect 449 1887 461 1921
rect 403 1853 461 1887
rect 403 1819 415 1853
rect 449 1819 461 1853
rect 403 1785 461 1819
rect 403 1751 415 1785
rect 449 1751 461 1785
rect 403 1717 461 1751
rect 403 1683 415 1717
rect 449 1683 461 1717
rect 403 1649 461 1683
rect 403 1615 415 1649
rect 449 1615 461 1649
rect 403 1581 461 1615
rect 403 1547 415 1581
rect 449 1547 461 1581
rect 403 1513 461 1547
rect 403 1479 415 1513
rect 449 1479 461 1513
rect 403 1445 461 1479
rect 403 1411 415 1445
rect 449 1411 461 1445
rect 403 1377 461 1411
rect 403 1343 415 1377
rect 449 1343 461 1377
rect 403 1309 461 1343
rect 403 1275 415 1309
rect 449 1275 461 1309
rect 403 1241 461 1275
rect 403 1207 415 1241
rect 449 1207 461 1241
rect 403 1173 461 1207
rect 403 1139 415 1173
rect 449 1139 461 1173
rect 403 1105 461 1139
rect 403 1071 415 1105
rect 449 1071 461 1105
rect 403 1037 461 1071
rect 403 1003 415 1037
rect 449 1003 461 1037
rect 403 969 461 1003
rect 403 935 415 969
rect 449 935 461 969
rect 403 901 461 935
rect 403 867 415 901
rect 449 867 461 901
rect 403 833 461 867
rect 403 799 415 833
rect 449 799 461 833
rect 403 765 461 799
rect 403 731 415 765
rect 449 731 461 765
rect 403 697 461 731
rect 403 663 415 697
rect 449 663 461 697
rect 403 629 461 663
rect 403 595 415 629
rect 449 595 461 629
rect 403 561 461 595
rect 403 527 415 561
rect 449 527 461 561
rect 403 493 461 527
rect 403 459 415 493
rect 449 459 461 493
rect 403 425 461 459
rect 403 391 415 425
rect 449 391 461 425
rect 403 357 461 391
rect 403 323 415 357
rect 449 323 461 357
rect 403 289 461 323
rect 403 255 415 289
rect 449 255 461 289
rect 403 221 461 255
rect 403 187 415 221
rect 449 187 461 221
rect 403 153 461 187
rect 403 119 415 153
rect 449 119 461 153
rect 403 85 461 119
rect 403 51 415 85
rect 449 51 461 85
rect 403 17 461 51
rect 403 -17 415 17
rect 449 -17 461 17
rect 403 -51 461 -17
rect 403 -85 415 -51
rect 449 -85 461 -51
rect 403 -119 461 -85
rect 403 -153 415 -119
rect 449 -153 461 -119
rect 403 -187 461 -153
rect 403 -221 415 -187
rect 449 -221 461 -187
rect 403 -255 461 -221
rect 403 -289 415 -255
rect 449 -289 461 -255
rect 403 -323 461 -289
rect 403 -357 415 -323
rect 449 -357 461 -323
rect 403 -391 461 -357
rect 403 -425 415 -391
rect 449 -425 461 -391
rect 403 -459 461 -425
rect 403 -493 415 -459
rect 449 -493 461 -459
rect 403 -527 461 -493
rect 403 -561 415 -527
rect 449 -561 461 -527
rect 403 -595 461 -561
rect 403 -629 415 -595
rect 449 -629 461 -595
rect 403 -663 461 -629
rect 403 -697 415 -663
rect 449 -697 461 -663
rect 403 -731 461 -697
rect 403 -765 415 -731
rect 449 -765 461 -731
rect 403 -799 461 -765
rect 403 -833 415 -799
rect 449 -833 461 -799
rect 403 -867 461 -833
rect 403 -901 415 -867
rect 449 -901 461 -867
rect 403 -935 461 -901
rect 403 -969 415 -935
rect 449 -969 461 -935
rect 403 -1003 461 -969
rect 403 -1037 415 -1003
rect 449 -1037 461 -1003
rect 403 -1071 461 -1037
rect 403 -1105 415 -1071
rect 449 -1105 461 -1071
rect 403 -1139 461 -1105
rect 403 -1173 415 -1139
rect 449 -1173 461 -1139
rect 403 -1207 461 -1173
rect 403 -1241 415 -1207
rect 449 -1241 461 -1207
rect 403 -1275 461 -1241
rect 403 -1309 415 -1275
rect 449 -1309 461 -1275
rect 403 -1343 461 -1309
rect 403 -1377 415 -1343
rect 449 -1377 461 -1343
rect 403 -1411 461 -1377
rect 403 -1445 415 -1411
rect 449 -1445 461 -1411
rect 403 -1479 461 -1445
rect 403 -1513 415 -1479
rect 449 -1513 461 -1479
rect 403 -1547 461 -1513
rect 403 -1581 415 -1547
rect 449 -1581 461 -1547
rect 403 -1615 461 -1581
rect 403 -1649 415 -1615
rect 449 -1649 461 -1615
rect 403 -1683 461 -1649
rect 403 -1717 415 -1683
rect 449 -1717 461 -1683
rect 403 -1751 461 -1717
rect 403 -1785 415 -1751
rect 449 -1785 461 -1751
rect 403 -1819 461 -1785
rect 403 -1853 415 -1819
rect 449 -1853 461 -1819
rect 403 -1887 461 -1853
rect 403 -1921 415 -1887
rect 449 -1921 461 -1887
rect 403 -1955 461 -1921
rect 403 -1989 415 -1955
rect 449 -1989 461 -1955
rect 403 -2023 461 -1989
rect 403 -2057 415 -2023
rect 449 -2057 461 -2023
rect 403 -2091 461 -2057
rect 403 -2125 415 -2091
rect 449 -2125 461 -2091
rect 403 -2159 461 -2125
rect 403 -2193 415 -2159
rect 449 -2193 461 -2159
rect 403 -2227 461 -2193
rect 403 -2261 415 -2227
rect 449 -2261 461 -2227
rect 403 -2295 461 -2261
rect 403 -2329 415 -2295
rect 449 -2329 461 -2295
rect 403 -2363 461 -2329
rect 403 -2397 415 -2363
rect 449 -2397 461 -2363
rect 403 -2431 461 -2397
rect 403 -2465 415 -2431
rect 449 -2465 461 -2431
rect 403 -2500 461 -2465
<< pdiffc >>
rect -449 2431 -415 2465
rect -449 2363 -415 2397
rect -449 2295 -415 2329
rect -449 2227 -415 2261
rect -449 2159 -415 2193
rect -449 2091 -415 2125
rect -449 2023 -415 2057
rect -449 1955 -415 1989
rect -449 1887 -415 1921
rect -449 1819 -415 1853
rect -449 1751 -415 1785
rect -449 1683 -415 1717
rect -449 1615 -415 1649
rect -449 1547 -415 1581
rect -449 1479 -415 1513
rect -449 1411 -415 1445
rect -449 1343 -415 1377
rect -449 1275 -415 1309
rect -449 1207 -415 1241
rect -449 1139 -415 1173
rect -449 1071 -415 1105
rect -449 1003 -415 1037
rect -449 935 -415 969
rect -449 867 -415 901
rect -449 799 -415 833
rect -449 731 -415 765
rect -449 663 -415 697
rect -449 595 -415 629
rect -449 527 -415 561
rect -449 459 -415 493
rect -449 391 -415 425
rect -449 323 -415 357
rect -449 255 -415 289
rect -449 187 -415 221
rect -449 119 -415 153
rect -449 51 -415 85
rect -449 -17 -415 17
rect -449 -85 -415 -51
rect -449 -153 -415 -119
rect -449 -221 -415 -187
rect -449 -289 -415 -255
rect -449 -357 -415 -323
rect -449 -425 -415 -391
rect -449 -493 -415 -459
rect -449 -561 -415 -527
rect -449 -629 -415 -595
rect -449 -697 -415 -663
rect -449 -765 -415 -731
rect -449 -833 -415 -799
rect -449 -901 -415 -867
rect -449 -969 -415 -935
rect -449 -1037 -415 -1003
rect -449 -1105 -415 -1071
rect -449 -1173 -415 -1139
rect -449 -1241 -415 -1207
rect -449 -1309 -415 -1275
rect -449 -1377 -415 -1343
rect -449 -1445 -415 -1411
rect -449 -1513 -415 -1479
rect -449 -1581 -415 -1547
rect -449 -1649 -415 -1615
rect -449 -1717 -415 -1683
rect -449 -1785 -415 -1751
rect -449 -1853 -415 -1819
rect -449 -1921 -415 -1887
rect -449 -1989 -415 -1955
rect -449 -2057 -415 -2023
rect -449 -2125 -415 -2091
rect -449 -2193 -415 -2159
rect -449 -2261 -415 -2227
rect -449 -2329 -415 -2295
rect -449 -2397 -415 -2363
rect -449 -2465 -415 -2431
rect -341 2431 -307 2465
rect -341 2363 -307 2397
rect -341 2295 -307 2329
rect -341 2227 -307 2261
rect -341 2159 -307 2193
rect -341 2091 -307 2125
rect -341 2023 -307 2057
rect -341 1955 -307 1989
rect -341 1887 -307 1921
rect -341 1819 -307 1853
rect -341 1751 -307 1785
rect -341 1683 -307 1717
rect -341 1615 -307 1649
rect -341 1547 -307 1581
rect -341 1479 -307 1513
rect -341 1411 -307 1445
rect -341 1343 -307 1377
rect -341 1275 -307 1309
rect -341 1207 -307 1241
rect -341 1139 -307 1173
rect -341 1071 -307 1105
rect -341 1003 -307 1037
rect -341 935 -307 969
rect -341 867 -307 901
rect -341 799 -307 833
rect -341 731 -307 765
rect -341 663 -307 697
rect -341 595 -307 629
rect -341 527 -307 561
rect -341 459 -307 493
rect -341 391 -307 425
rect -341 323 -307 357
rect -341 255 -307 289
rect -341 187 -307 221
rect -341 119 -307 153
rect -341 51 -307 85
rect -341 -17 -307 17
rect -341 -85 -307 -51
rect -341 -153 -307 -119
rect -341 -221 -307 -187
rect -341 -289 -307 -255
rect -341 -357 -307 -323
rect -341 -425 -307 -391
rect -341 -493 -307 -459
rect -341 -561 -307 -527
rect -341 -629 -307 -595
rect -341 -697 -307 -663
rect -341 -765 -307 -731
rect -341 -833 -307 -799
rect -341 -901 -307 -867
rect -341 -969 -307 -935
rect -341 -1037 -307 -1003
rect -341 -1105 -307 -1071
rect -341 -1173 -307 -1139
rect -341 -1241 -307 -1207
rect -341 -1309 -307 -1275
rect -341 -1377 -307 -1343
rect -341 -1445 -307 -1411
rect -341 -1513 -307 -1479
rect -341 -1581 -307 -1547
rect -341 -1649 -307 -1615
rect -341 -1717 -307 -1683
rect -341 -1785 -307 -1751
rect -341 -1853 -307 -1819
rect -341 -1921 -307 -1887
rect -341 -1989 -307 -1955
rect -341 -2057 -307 -2023
rect -341 -2125 -307 -2091
rect -341 -2193 -307 -2159
rect -341 -2261 -307 -2227
rect -341 -2329 -307 -2295
rect -341 -2397 -307 -2363
rect -341 -2465 -307 -2431
rect -233 2431 -199 2465
rect -233 2363 -199 2397
rect -233 2295 -199 2329
rect -233 2227 -199 2261
rect -233 2159 -199 2193
rect -233 2091 -199 2125
rect -233 2023 -199 2057
rect -233 1955 -199 1989
rect -233 1887 -199 1921
rect -233 1819 -199 1853
rect -233 1751 -199 1785
rect -233 1683 -199 1717
rect -233 1615 -199 1649
rect -233 1547 -199 1581
rect -233 1479 -199 1513
rect -233 1411 -199 1445
rect -233 1343 -199 1377
rect -233 1275 -199 1309
rect -233 1207 -199 1241
rect -233 1139 -199 1173
rect -233 1071 -199 1105
rect -233 1003 -199 1037
rect -233 935 -199 969
rect -233 867 -199 901
rect -233 799 -199 833
rect -233 731 -199 765
rect -233 663 -199 697
rect -233 595 -199 629
rect -233 527 -199 561
rect -233 459 -199 493
rect -233 391 -199 425
rect -233 323 -199 357
rect -233 255 -199 289
rect -233 187 -199 221
rect -233 119 -199 153
rect -233 51 -199 85
rect -233 -17 -199 17
rect -233 -85 -199 -51
rect -233 -153 -199 -119
rect -233 -221 -199 -187
rect -233 -289 -199 -255
rect -233 -357 -199 -323
rect -233 -425 -199 -391
rect -233 -493 -199 -459
rect -233 -561 -199 -527
rect -233 -629 -199 -595
rect -233 -697 -199 -663
rect -233 -765 -199 -731
rect -233 -833 -199 -799
rect -233 -901 -199 -867
rect -233 -969 -199 -935
rect -233 -1037 -199 -1003
rect -233 -1105 -199 -1071
rect -233 -1173 -199 -1139
rect -233 -1241 -199 -1207
rect -233 -1309 -199 -1275
rect -233 -1377 -199 -1343
rect -233 -1445 -199 -1411
rect -233 -1513 -199 -1479
rect -233 -1581 -199 -1547
rect -233 -1649 -199 -1615
rect -233 -1717 -199 -1683
rect -233 -1785 -199 -1751
rect -233 -1853 -199 -1819
rect -233 -1921 -199 -1887
rect -233 -1989 -199 -1955
rect -233 -2057 -199 -2023
rect -233 -2125 -199 -2091
rect -233 -2193 -199 -2159
rect -233 -2261 -199 -2227
rect -233 -2329 -199 -2295
rect -233 -2397 -199 -2363
rect -233 -2465 -199 -2431
rect -125 2431 -91 2465
rect -125 2363 -91 2397
rect -125 2295 -91 2329
rect -125 2227 -91 2261
rect -125 2159 -91 2193
rect -125 2091 -91 2125
rect -125 2023 -91 2057
rect -125 1955 -91 1989
rect -125 1887 -91 1921
rect -125 1819 -91 1853
rect -125 1751 -91 1785
rect -125 1683 -91 1717
rect -125 1615 -91 1649
rect -125 1547 -91 1581
rect -125 1479 -91 1513
rect -125 1411 -91 1445
rect -125 1343 -91 1377
rect -125 1275 -91 1309
rect -125 1207 -91 1241
rect -125 1139 -91 1173
rect -125 1071 -91 1105
rect -125 1003 -91 1037
rect -125 935 -91 969
rect -125 867 -91 901
rect -125 799 -91 833
rect -125 731 -91 765
rect -125 663 -91 697
rect -125 595 -91 629
rect -125 527 -91 561
rect -125 459 -91 493
rect -125 391 -91 425
rect -125 323 -91 357
rect -125 255 -91 289
rect -125 187 -91 221
rect -125 119 -91 153
rect -125 51 -91 85
rect -125 -17 -91 17
rect -125 -85 -91 -51
rect -125 -153 -91 -119
rect -125 -221 -91 -187
rect -125 -289 -91 -255
rect -125 -357 -91 -323
rect -125 -425 -91 -391
rect -125 -493 -91 -459
rect -125 -561 -91 -527
rect -125 -629 -91 -595
rect -125 -697 -91 -663
rect -125 -765 -91 -731
rect -125 -833 -91 -799
rect -125 -901 -91 -867
rect -125 -969 -91 -935
rect -125 -1037 -91 -1003
rect -125 -1105 -91 -1071
rect -125 -1173 -91 -1139
rect -125 -1241 -91 -1207
rect -125 -1309 -91 -1275
rect -125 -1377 -91 -1343
rect -125 -1445 -91 -1411
rect -125 -1513 -91 -1479
rect -125 -1581 -91 -1547
rect -125 -1649 -91 -1615
rect -125 -1717 -91 -1683
rect -125 -1785 -91 -1751
rect -125 -1853 -91 -1819
rect -125 -1921 -91 -1887
rect -125 -1989 -91 -1955
rect -125 -2057 -91 -2023
rect -125 -2125 -91 -2091
rect -125 -2193 -91 -2159
rect -125 -2261 -91 -2227
rect -125 -2329 -91 -2295
rect -125 -2397 -91 -2363
rect -125 -2465 -91 -2431
rect -17 2431 17 2465
rect -17 2363 17 2397
rect -17 2295 17 2329
rect -17 2227 17 2261
rect -17 2159 17 2193
rect -17 2091 17 2125
rect -17 2023 17 2057
rect -17 1955 17 1989
rect -17 1887 17 1921
rect -17 1819 17 1853
rect -17 1751 17 1785
rect -17 1683 17 1717
rect -17 1615 17 1649
rect -17 1547 17 1581
rect -17 1479 17 1513
rect -17 1411 17 1445
rect -17 1343 17 1377
rect -17 1275 17 1309
rect -17 1207 17 1241
rect -17 1139 17 1173
rect -17 1071 17 1105
rect -17 1003 17 1037
rect -17 935 17 969
rect -17 867 17 901
rect -17 799 17 833
rect -17 731 17 765
rect -17 663 17 697
rect -17 595 17 629
rect -17 527 17 561
rect -17 459 17 493
rect -17 391 17 425
rect -17 323 17 357
rect -17 255 17 289
rect -17 187 17 221
rect -17 119 17 153
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect -17 -153 17 -119
rect -17 -221 17 -187
rect -17 -289 17 -255
rect -17 -357 17 -323
rect -17 -425 17 -391
rect -17 -493 17 -459
rect -17 -561 17 -527
rect -17 -629 17 -595
rect -17 -697 17 -663
rect -17 -765 17 -731
rect -17 -833 17 -799
rect -17 -901 17 -867
rect -17 -969 17 -935
rect -17 -1037 17 -1003
rect -17 -1105 17 -1071
rect -17 -1173 17 -1139
rect -17 -1241 17 -1207
rect -17 -1309 17 -1275
rect -17 -1377 17 -1343
rect -17 -1445 17 -1411
rect -17 -1513 17 -1479
rect -17 -1581 17 -1547
rect -17 -1649 17 -1615
rect -17 -1717 17 -1683
rect -17 -1785 17 -1751
rect -17 -1853 17 -1819
rect -17 -1921 17 -1887
rect -17 -1989 17 -1955
rect -17 -2057 17 -2023
rect -17 -2125 17 -2091
rect -17 -2193 17 -2159
rect -17 -2261 17 -2227
rect -17 -2329 17 -2295
rect -17 -2397 17 -2363
rect -17 -2465 17 -2431
rect 91 2431 125 2465
rect 91 2363 125 2397
rect 91 2295 125 2329
rect 91 2227 125 2261
rect 91 2159 125 2193
rect 91 2091 125 2125
rect 91 2023 125 2057
rect 91 1955 125 1989
rect 91 1887 125 1921
rect 91 1819 125 1853
rect 91 1751 125 1785
rect 91 1683 125 1717
rect 91 1615 125 1649
rect 91 1547 125 1581
rect 91 1479 125 1513
rect 91 1411 125 1445
rect 91 1343 125 1377
rect 91 1275 125 1309
rect 91 1207 125 1241
rect 91 1139 125 1173
rect 91 1071 125 1105
rect 91 1003 125 1037
rect 91 935 125 969
rect 91 867 125 901
rect 91 799 125 833
rect 91 731 125 765
rect 91 663 125 697
rect 91 595 125 629
rect 91 527 125 561
rect 91 459 125 493
rect 91 391 125 425
rect 91 323 125 357
rect 91 255 125 289
rect 91 187 125 221
rect 91 119 125 153
rect 91 51 125 85
rect 91 -17 125 17
rect 91 -85 125 -51
rect 91 -153 125 -119
rect 91 -221 125 -187
rect 91 -289 125 -255
rect 91 -357 125 -323
rect 91 -425 125 -391
rect 91 -493 125 -459
rect 91 -561 125 -527
rect 91 -629 125 -595
rect 91 -697 125 -663
rect 91 -765 125 -731
rect 91 -833 125 -799
rect 91 -901 125 -867
rect 91 -969 125 -935
rect 91 -1037 125 -1003
rect 91 -1105 125 -1071
rect 91 -1173 125 -1139
rect 91 -1241 125 -1207
rect 91 -1309 125 -1275
rect 91 -1377 125 -1343
rect 91 -1445 125 -1411
rect 91 -1513 125 -1479
rect 91 -1581 125 -1547
rect 91 -1649 125 -1615
rect 91 -1717 125 -1683
rect 91 -1785 125 -1751
rect 91 -1853 125 -1819
rect 91 -1921 125 -1887
rect 91 -1989 125 -1955
rect 91 -2057 125 -2023
rect 91 -2125 125 -2091
rect 91 -2193 125 -2159
rect 91 -2261 125 -2227
rect 91 -2329 125 -2295
rect 91 -2397 125 -2363
rect 91 -2465 125 -2431
rect 199 2431 233 2465
rect 199 2363 233 2397
rect 199 2295 233 2329
rect 199 2227 233 2261
rect 199 2159 233 2193
rect 199 2091 233 2125
rect 199 2023 233 2057
rect 199 1955 233 1989
rect 199 1887 233 1921
rect 199 1819 233 1853
rect 199 1751 233 1785
rect 199 1683 233 1717
rect 199 1615 233 1649
rect 199 1547 233 1581
rect 199 1479 233 1513
rect 199 1411 233 1445
rect 199 1343 233 1377
rect 199 1275 233 1309
rect 199 1207 233 1241
rect 199 1139 233 1173
rect 199 1071 233 1105
rect 199 1003 233 1037
rect 199 935 233 969
rect 199 867 233 901
rect 199 799 233 833
rect 199 731 233 765
rect 199 663 233 697
rect 199 595 233 629
rect 199 527 233 561
rect 199 459 233 493
rect 199 391 233 425
rect 199 323 233 357
rect 199 255 233 289
rect 199 187 233 221
rect 199 119 233 153
rect 199 51 233 85
rect 199 -17 233 17
rect 199 -85 233 -51
rect 199 -153 233 -119
rect 199 -221 233 -187
rect 199 -289 233 -255
rect 199 -357 233 -323
rect 199 -425 233 -391
rect 199 -493 233 -459
rect 199 -561 233 -527
rect 199 -629 233 -595
rect 199 -697 233 -663
rect 199 -765 233 -731
rect 199 -833 233 -799
rect 199 -901 233 -867
rect 199 -969 233 -935
rect 199 -1037 233 -1003
rect 199 -1105 233 -1071
rect 199 -1173 233 -1139
rect 199 -1241 233 -1207
rect 199 -1309 233 -1275
rect 199 -1377 233 -1343
rect 199 -1445 233 -1411
rect 199 -1513 233 -1479
rect 199 -1581 233 -1547
rect 199 -1649 233 -1615
rect 199 -1717 233 -1683
rect 199 -1785 233 -1751
rect 199 -1853 233 -1819
rect 199 -1921 233 -1887
rect 199 -1989 233 -1955
rect 199 -2057 233 -2023
rect 199 -2125 233 -2091
rect 199 -2193 233 -2159
rect 199 -2261 233 -2227
rect 199 -2329 233 -2295
rect 199 -2397 233 -2363
rect 199 -2465 233 -2431
rect 307 2431 341 2465
rect 307 2363 341 2397
rect 307 2295 341 2329
rect 307 2227 341 2261
rect 307 2159 341 2193
rect 307 2091 341 2125
rect 307 2023 341 2057
rect 307 1955 341 1989
rect 307 1887 341 1921
rect 307 1819 341 1853
rect 307 1751 341 1785
rect 307 1683 341 1717
rect 307 1615 341 1649
rect 307 1547 341 1581
rect 307 1479 341 1513
rect 307 1411 341 1445
rect 307 1343 341 1377
rect 307 1275 341 1309
rect 307 1207 341 1241
rect 307 1139 341 1173
rect 307 1071 341 1105
rect 307 1003 341 1037
rect 307 935 341 969
rect 307 867 341 901
rect 307 799 341 833
rect 307 731 341 765
rect 307 663 341 697
rect 307 595 341 629
rect 307 527 341 561
rect 307 459 341 493
rect 307 391 341 425
rect 307 323 341 357
rect 307 255 341 289
rect 307 187 341 221
rect 307 119 341 153
rect 307 51 341 85
rect 307 -17 341 17
rect 307 -85 341 -51
rect 307 -153 341 -119
rect 307 -221 341 -187
rect 307 -289 341 -255
rect 307 -357 341 -323
rect 307 -425 341 -391
rect 307 -493 341 -459
rect 307 -561 341 -527
rect 307 -629 341 -595
rect 307 -697 341 -663
rect 307 -765 341 -731
rect 307 -833 341 -799
rect 307 -901 341 -867
rect 307 -969 341 -935
rect 307 -1037 341 -1003
rect 307 -1105 341 -1071
rect 307 -1173 341 -1139
rect 307 -1241 341 -1207
rect 307 -1309 341 -1275
rect 307 -1377 341 -1343
rect 307 -1445 341 -1411
rect 307 -1513 341 -1479
rect 307 -1581 341 -1547
rect 307 -1649 341 -1615
rect 307 -1717 341 -1683
rect 307 -1785 341 -1751
rect 307 -1853 341 -1819
rect 307 -1921 341 -1887
rect 307 -1989 341 -1955
rect 307 -2057 341 -2023
rect 307 -2125 341 -2091
rect 307 -2193 341 -2159
rect 307 -2261 341 -2227
rect 307 -2329 341 -2295
rect 307 -2397 341 -2363
rect 307 -2465 341 -2431
rect 415 2431 449 2465
rect 415 2363 449 2397
rect 415 2295 449 2329
rect 415 2227 449 2261
rect 415 2159 449 2193
rect 415 2091 449 2125
rect 415 2023 449 2057
rect 415 1955 449 1989
rect 415 1887 449 1921
rect 415 1819 449 1853
rect 415 1751 449 1785
rect 415 1683 449 1717
rect 415 1615 449 1649
rect 415 1547 449 1581
rect 415 1479 449 1513
rect 415 1411 449 1445
rect 415 1343 449 1377
rect 415 1275 449 1309
rect 415 1207 449 1241
rect 415 1139 449 1173
rect 415 1071 449 1105
rect 415 1003 449 1037
rect 415 935 449 969
rect 415 867 449 901
rect 415 799 449 833
rect 415 731 449 765
rect 415 663 449 697
rect 415 595 449 629
rect 415 527 449 561
rect 415 459 449 493
rect 415 391 449 425
rect 415 323 449 357
rect 415 255 449 289
rect 415 187 449 221
rect 415 119 449 153
rect 415 51 449 85
rect 415 -17 449 17
rect 415 -85 449 -51
rect 415 -153 449 -119
rect 415 -221 449 -187
rect 415 -289 449 -255
rect 415 -357 449 -323
rect 415 -425 449 -391
rect 415 -493 449 -459
rect 415 -561 449 -527
rect 415 -629 449 -595
rect 415 -697 449 -663
rect 415 -765 449 -731
rect 415 -833 449 -799
rect 415 -901 449 -867
rect 415 -969 449 -935
rect 415 -1037 449 -1003
rect 415 -1105 449 -1071
rect 415 -1173 449 -1139
rect 415 -1241 449 -1207
rect 415 -1309 449 -1275
rect 415 -1377 449 -1343
rect 415 -1445 449 -1411
rect 415 -1513 449 -1479
rect 415 -1581 449 -1547
rect 415 -1649 449 -1615
rect 415 -1717 449 -1683
rect 415 -1785 449 -1751
rect 415 -1853 449 -1819
rect 415 -1921 449 -1887
rect 415 -1989 449 -1955
rect 415 -2057 449 -2023
rect 415 -2125 449 -2091
rect 415 -2193 449 -2159
rect 415 -2261 449 -2227
rect 415 -2329 449 -2295
rect 415 -2397 449 -2363
rect 415 -2465 449 -2431
<< nsubdiff >>
rect -563 2649 -459 2683
rect -425 2649 -391 2683
rect -357 2649 -323 2683
rect -289 2649 -255 2683
rect -221 2649 -187 2683
rect -153 2649 -119 2683
rect -85 2649 -51 2683
rect -17 2649 17 2683
rect 51 2649 85 2683
rect 119 2649 153 2683
rect 187 2649 221 2683
rect 255 2649 289 2683
rect 323 2649 357 2683
rect 391 2649 425 2683
rect 459 2649 563 2683
rect -563 2567 -529 2649
rect -563 2499 -529 2533
rect 529 2567 563 2649
rect -563 2431 -529 2465
rect -563 2363 -529 2397
rect -563 2295 -529 2329
rect -563 2227 -529 2261
rect -563 2159 -529 2193
rect -563 2091 -529 2125
rect -563 2023 -529 2057
rect -563 1955 -529 1989
rect -563 1887 -529 1921
rect -563 1819 -529 1853
rect -563 1751 -529 1785
rect -563 1683 -529 1717
rect -563 1615 -529 1649
rect -563 1547 -529 1581
rect -563 1479 -529 1513
rect -563 1411 -529 1445
rect -563 1343 -529 1377
rect -563 1275 -529 1309
rect -563 1207 -529 1241
rect -563 1139 -529 1173
rect -563 1071 -529 1105
rect -563 1003 -529 1037
rect -563 935 -529 969
rect -563 867 -529 901
rect -563 799 -529 833
rect -563 731 -529 765
rect -563 663 -529 697
rect -563 595 -529 629
rect -563 527 -529 561
rect -563 459 -529 493
rect -563 391 -529 425
rect -563 323 -529 357
rect -563 255 -529 289
rect -563 187 -529 221
rect -563 119 -529 153
rect -563 51 -529 85
rect -563 -17 -529 17
rect -563 -85 -529 -51
rect -563 -153 -529 -119
rect -563 -221 -529 -187
rect -563 -289 -529 -255
rect -563 -357 -529 -323
rect -563 -425 -529 -391
rect -563 -493 -529 -459
rect -563 -561 -529 -527
rect -563 -629 -529 -595
rect -563 -697 -529 -663
rect -563 -765 -529 -731
rect -563 -833 -529 -799
rect -563 -901 -529 -867
rect -563 -969 -529 -935
rect -563 -1037 -529 -1003
rect -563 -1105 -529 -1071
rect -563 -1173 -529 -1139
rect -563 -1241 -529 -1207
rect -563 -1309 -529 -1275
rect -563 -1377 -529 -1343
rect -563 -1445 -529 -1411
rect -563 -1513 -529 -1479
rect -563 -1581 -529 -1547
rect -563 -1649 -529 -1615
rect -563 -1717 -529 -1683
rect -563 -1785 -529 -1751
rect -563 -1853 -529 -1819
rect -563 -1921 -529 -1887
rect -563 -1989 -529 -1955
rect -563 -2057 -529 -2023
rect -563 -2125 -529 -2091
rect -563 -2193 -529 -2159
rect -563 -2261 -529 -2227
rect -563 -2329 -529 -2295
rect -563 -2397 -529 -2363
rect -563 -2465 -529 -2431
rect -563 -2533 -529 -2499
rect 529 2499 563 2533
rect 529 2431 563 2465
rect 529 2363 563 2397
rect 529 2295 563 2329
rect 529 2227 563 2261
rect 529 2159 563 2193
rect 529 2091 563 2125
rect 529 2023 563 2057
rect 529 1955 563 1989
rect 529 1887 563 1921
rect 529 1819 563 1853
rect 529 1751 563 1785
rect 529 1683 563 1717
rect 529 1615 563 1649
rect 529 1547 563 1581
rect 529 1479 563 1513
rect 529 1411 563 1445
rect 529 1343 563 1377
rect 529 1275 563 1309
rect 529 1207 563 1241
rect 529 1139 563 1173
rect 529 1071 563 1105
rect 529 1003 563 1037
rect 529 935 563 969
rect 529 867 563 901
rect 529 799 563 833
rect 529 731 563 765
rect 529 663 563 697
rect 529 595 563 629
rect 529 527 563 561
rect 529 459 563 493
rect 529 391 563 425
rect 529 323 563 357
rect 529 255 563 289
rect 529 187 563 221
rect 529 119 563 153
rect 529 51 563 85
rect 529 -17 563 17
rect 529 -85 563 -51
rect 529 -153 563 -119
rect 529 -221 563 -187
rect 529 -289 563 -255
rect 529 -357 563 -323
rect 529 -425 563 -391
rect 529 -493 563 -459
rect 529 -561 563 -527
rect 529 -629 563 -595
rect 529 -697 563 -663
rect 529 -765 563 -731
rect 529 -833 563 -799
rect 529 -901 563 -867
rect 529 -969 563 -935
rect 529 -1037 563 -1003
rect 529 -1105 563 -1071
rect 529 -1173 563 -1139
rect 529 -1241 563 -1207
rect 529 -1309 563 -1275
rect 529 -1377 563 -1343
rect 529 -1445 563 -1411
rect 529 -1513 563 -1479
rect 529 -1581 563 -1547
rect 529 -1649 563 -1615
rect 529 -1717 563 -1683
rect 529 -1785 563 -1751
rect 529 -1853 563 -1819
rect 529 -1921 563 -1887
rect 529 -1989 563 -1955
rect 529 -2057 563 -2023
rect 529 -2125 563 -2091
rect 529 -2193 563 -2159
rect 529 -2261 563 -2227
rect 529 -2329 563 -2295
rect 529 -2397 563 -2363
rect 529 -2465 563 -2431
rect -563 -2649 -529 -2567
rect 529 -2533 563 -2499
rect 529 -2649 563 -2567
rect -563 -2683 -459 -2649
rect -425 -2683 -391 -2649
rect -357 -2683 -323 -2649
rect -289 -2683 -255 -2649
rect -221 -2683 -187 -2649
rect -153 -2683 -119 -2649
rect -85 -2683 -51 -2649
rect -17 -2683 17 -2649
rect 51 -2683 85 -2649
rect 119 -2683 153 -2649
rect 187 -2683 221 -2649
rect 255 -2683 289 -2649
rect 323 -2683 357 -2649
rect 391 -2683 425 -2649
rect 459 -2683 563 -2649
<< nsubdiffcont >>
rect -459 2649 -425 2683
rect -391 2649 -357 2683
rect -323 2649 -289 2683
rect -255 2649 -221 2683
rect -187 2649 -153 2683
rect -119 2649 -85 2683
rect -51 2649 -17 2683
rect 17 2649 51 2683
rect 85 2649 119 2683
rect 153 2649 187 2683
rect 221 2649 255 2683
rect 289 2649 323 2683
rect 357 2649 391 2683
rect 425 2649 459 2683
rect -563 2533 -529 2567
rect 529 2533 563 2567
rect -563 2465 -529 2499
rect -563 2397 -529 2431
rect -563 2329 -529 2363
rect -563 2261 -529 2295
rect -563 2193 -529 2227
rect -563 2125 -529 2159
rect -563 2057 -529 2091
rect -563 1989 -529 2023
rect -563 1921 -529 1955
rect -563 1853 -529 1887
rect -563 1785 -529 1819
rect -563 1717 -529 1751
rect -563 1649 -529 1683
rect -563 1581 -529 1615
rect -563 1513 -529 1547
rect -563 1445 -529 1479
rect -563 1377 -529 1411
rect -563 1309 -529 1343
rect -563 1241 -529 1275
rect -563 1173 -529 1207
rect -563 1105 -529 1139
rect -563 1037 -529 1071
rect -563 969 -529 1003
rect -563 901 -529 935
rect -563 833 -529 867
rect -563 765 -529 799
rect -563 697 -529 731
rect -563 629 -529 663
rect -563 561 -529 595
rect -563 493 -529 527
rect -563 425 -529 459
rect -563 357 -529 391
rect -563 289 -529 323
rect -563 221 -529 255
rect -563 153 -529 187
rect -563 85 -529 119
rect -563 17 -529 51
rect -563 -51 -529 -17
rect -563 -119 -529 -85
rect -563 -187 -529 -153
rect -563 -255 -529 -221
rect -563 -323 -529 -289
rect -563 -391 -529 -357
rect -563 -459 -529 -425
rect -563 -527 -529 -493
rect -563 -595 -529 -561
rect -563 -663 -529 -629
rect -563 -731 -529 -697
rect -563 -799 -529 -765
rect -563 -867 -529 -833
rect -563 -935 -529 -901
rect -563 -1003 -529 -969
rect -563 -1071 -529 -1037
rect -563 -1139 -529 -1105
rect -563 -1207 -529 -1173
rect -563 -1275 -529 -1241
rect -563 -1343 -529 -1309
rect -563 -1411 -529 -1377
rect -563 -1479 -529 -1445
rect -563 -1547 -529 -1513
rect -563 -1615 -529 -1581
rect -563 -1683 -529 -1649
rect -563 -1751 -529 -1717
rect -563 -1819 -529 -1785
rect -563 -1887 -529 -1853
rect -563 -1955 -529 -1921
rect -563 -2023 -529 -1989
rect -563 -2091 -529 -2057
rect -563 -2159 -529 -2125
rect -563 -2227 -529 -2193
rect -563 -2295 -529 -2261
rect -563 -2363 -529 -2329
rect -563 -2431 -529 -2397
rect -563 -2499 -529 -2465
rect 529 2465 563 2499
rect 529 2397 563 2431
rect 529 2329 563 2363
rect 529 2261 563 2295
rect 529 2193 563 2227
rect 529 2125 563 2159
rect 529 2057 563 2091
rect 529 1989 563 2023
rect 529 1921 563 1955
rect 529 1853 563 1887
rect 529 1785 563 1819
rect 529 1717 563 1751
rect 529 1649 563 1683
rect 529 1581 563 1615
rect 529 1513 563 1547
rect 529 1445 563 1479
rect 529 1377 563 1411
rect 529 1309 563 1343
rect 529 1241 563 1275
rect 529 1173 563 1207
rect 529 1105 563 1139
rect 529 1037 563 1071
rect 529 969 563 1003
rect 529 901 563 935
rect 529 833 563 867
rect 529 765 563 799
rect 529 697 563 731
rect 529 629 563 663
rect 529 561 563 595
rect 529 493 563 527
rect 529 425 563 459
rect 529 357 563 391
rect 529 289 563 323
rect 529 221 563 255
rect 529 153 563 187
rect 529 85 563 119
rect 529 17 563 51
rect 529 -51 563 -17
rect 529 -119 563 -85
rect 529 -187 563 -153
rect 529 -255 563 -221
rect 529 -323 563 -289
rect 529 -391 563 -357
rect 529 -459 563 -425
rect 529 -527 563 -493
rect 529 -595 563 -561
rect 529 -663 563 -629
rect 529 -731 563 -697
rect 529 -799 563 -765
rect 529 -867 563 -833
rect 529 -935 563 -901
rect 529 -1003 563 -969
rect 529 -1071 563 -1037
rect 529 -1139 563 -1105
rect 529 -1207 563 -1173
rect 529 -1275 563 -1241
rect 529 -1343 563 -1309
rect 529 -1411 563 -1377
rect 529 -1479 563 -1445
rect 529 -1547 563 -1513
rect 529 -1615 563 -1581
rect 529 -1683 563 -1649
rect 529 -1751 563 -1717
rect 529 -1819 563 -1785
rect 529 -1887 563 -1853
rect 529 -1955 563 -1921
rect 529 -2023 563 -1989
rect 529 -2091 563 -2057
rect 529 -2159 563 -2125
rect 529 -2227 563 -2193
rect 529 -2295 563 -2261
rect 529 -2363 563 -2329
rect 529 -2431 563 -2397
rect 529 -2499 563 -2465
rect -563 -2567 -529 -2533
rect 529 -2567 563 -2533
rect -459 -2683 -425 -2649
rect -391 -2683 -357 -2649
rect -323 -2683 -289 -2649
rect -255 -2683 -221 -2649
rect -187 -2683 -153 -2649
rect -119 -2683 -85 -2649
rect -51 -2683 -17 -2649
rect 17 -2683 51 -2649
rect 85 -2683 119 -2649
rect 153 -2683 187 -2649
rect 221 -2683 255 -2649
rect 289 -2683 323 -2649
rect 357 -2683 391 -2649
rect 425 -2683 459 -2649
<< poly >>
rect -303 2581 -237 2597
rect -303 2547 -287 2581
rect -253 2547 -237 2581
rect -303 2531 -237 2547
rect -87 2581 -21 2597
rect -87 2547 -71 2581
rect -37 2547 -21 2581
rect -87 2531 -21 2547
rect 129 2581 195 2597
rect 129 2547 145 2581
rect 179 2547 195 2581
rect 129 2531 195 2547
rect 345 2581 411 2597
rect 345 2547 361 2581
rect 395 2547 411 2581
rect 345 2531 411 2547
rect -403 2500 -353 2526
rect -295 2500 -245 2531
rect -187 2500 -137 2526
rect -79 2500 -29 2531
rect 29 2500 79 2526
rect 137 2500 187 2531
rect 245 2500 295 2526
rect 353 2500 403 2531
rect -403 -2531 -353 -2500
rect -295 -2526 -245 -2500
rect -187 -2531 -137 -2500
rect -79 -2526 -29 -2500
rect 29 -2531 79 -2500
rect 137 -2526 187 -2500
rect 245 -2531 295 -2500
rect 353 -2526 403 -2500
rect -411 -2547 -345 -2531
rect -411 -2581 -395 -2547
rect -361 -2581 -345 -2547
rect -411 -2597 -345 -2581
rect -195 -2547 -129 -2531
rect -195 -2581 -179 -2547
rect -145 -2581 -129 -2547
rect -195 -2597 -129 -2581
rect 21 -2547 87 -2531
rect 21 -2581 37 -2547
rect 71 -2581 87 -2547
rect 21 -2597 87 -2581
rect 237 -2547 303 -2531
rect 237 -2581 253 -2547
rect 287 -2581 303 -2547
rect 237 -2597 303 -2581
<< polycont >>
rect -287 2547 -253 2581
rect -71 2547 -37 2581
rect 145 2547 179 2581
rect 361 2547 395 2581
rect -395 -2581 -361 -2547
rect -179 -2581 -145 -2547
rect 37 -2581 71 -2547
rect 253 -2581 287 -2547
<< locali >>
rect -563 2649 -459 2683
rect -425 2649 -391 2683
rect -357 2649 -323 2683
rect -289 2649 -255 2683
rect -221 2649 -187 2683
rect -153 2649 -119 2683
rect -85 2649 -51 2683
rect -17 2649 17 2683
rect 51 2649 85 2683
rect 119 2649 153 2683
rect 187 2649 221 2683
rect 255 2649 289 2683
rect 323 2649 357 2683
rect 391 2649 425 2683
rect 459 2649 563 2683
rect -563 2567 -529 2649
rect -303 2547 -287 2581
rect -253 2547 -237 2581
rect -87 2547 -71 2581
rect -37 2547 -21 2581
rect 129 2547 145 2581
rect 179 2547 195 2581
rect 345 2547 361 2581
rect 395 2547 411 2581
rect 529 2567 563 2649
rect -563 2499 -529 2533
rect -563 2431 -529 2465
rect -563 2363 -529 2397
rect -563 2295 -529 2329
rect -563 2227 -529 2261
rect -563 2159 -529 2193
rect -563 2091 -529 2125
rect -563 2023 -529 2057
rect -563 1955 -529 1989
rect -563 1887 -529 1921
rect -563 1819 -529 1853
rect -563 1751 -529 1785
rect -563 1683 -529 1717
rect -563 1615 -529 1649
rect -563 1547 -529 1581
rect -563 1479 -529 1513
rect -563 1411 -529 1445
rect -563 1343 -529 1377
rect -563 1275 -529 1309
rect -563 1207 -529 1241
rect -563 1139 -529 1173
rect -563 1071 -529 1105
rect -563 1003 -529 1037
rect -563 935 -529 969
rect -563 867 -529 901
rect -563 799 -529 833
rect -563 731 -529 765
rect -563 663 -529 697
rect -563 595 -529 629
rect -563 527 -529 561
rect -563 459 -529 493
rect -563 391 -529 425
rect -563 323 -529 357
rect -563 255 -529 289
rect -563 187 -529 221
rect -563 119 -529 153
rect -563 51 -529 85
rect -563 -17 -529 17
rect -563 -85 -529 -51
rect -563 -153 -529 -119
rect -563 -221 -529 -187
rect -563 -289 -529 -255
rect -563 -357 -529 -323
rect -563 -425 -529 -391
rect -563 -493 -529 -459
rect -563 -561 -529 -527
rect -563 -629 -529 -595
rect -563 -697 -529 -663
rect -563 -765 -529 -731
rect -563 -833 -529 -799
rect -563 -901 -529 -867
rect -563 -969 -529 -935
rect -563 -1037 -529 -1003
rect -563 -1105 -529 -1071
rect -563 -1173 -529 -1139
rect -563 -1241 -529 -1207
rect -563 -1309 -529 -1275
rect -563 -1377 -529 -1343
rect -563 -1445 -529 -1411
rect -563 -1513 -529 -1479
rect -563 -1581 -529 -1547
rect -563 -1649 -529 -1615
rect -563 -1717 -529 -1683
rect -563 -1785 -529 -1751
rect -563 -1853 -529 -1819
rect -563 -1921 -529 -1887
rect -563 -1989 -529 -1955
rect -563 -2057 -529 -2023
rect -563 -2125 -529 -2091
rect -563 -2193 -529 -2159
rect -563 -2261 -529 -2227
rect -563 -2329 -529 -2295
rect -563 -2397 -529 -2363
rect -563 -2465 -529 -2431
rect -563 -2533 -529 -2499
rect -449 2465 -415 2504
rect -449 2397 -415 2431
rect -449 2329 -415 2359
rect -449 2261 -415 2287
rect -449 2193 -415 2215
rect -449 2125 -415 2143
rect -449 2057 -415 2071
rect -449 1989 -415 1999
rect -449 1921 -415 1927
rect -449 1853 -415 1855
rect -449 1817 -415 1819
rect -449 1745 -415 1751
rect -449 1673 -415 1683
rect -449 1601 -415 1615
rect -449 1529 -415 1547
rect -449 1457 -415 1479
rect -449 1385 -415 1411
rect -449 1313 -415 1343
rect -449 1241 -415 1275
rect -449 1173 -415 1207
rect -449 1105 -415 1135
rect -449 1037 -415 1063
rect -449 969 -415 991
rect -449 901 -415 919
rect -449 833 -415 847
rect -449 765 -415 775
rect -449 697 -415 703
rect -449 629 -415 631
rect -449 593 -415 595
rect -449 521 -415 527
rect -449 449 -415 459
rect -449 377 -415 391
rect -449 305 -415 323
rect -449 233 -415 255
rect -449 161 -415 187
rect -449 89 -415 119
rect -449 17 -415 51
rect -449 -51 -415 -17
rect -449 -119 -415 -89
rect -449 -187 -415 -161
rect -449 -255 -415 -233
rect -449 -323 -415 -305
rect -449 -391 -415 -377
rect -449 -459 -415 -449
rect -449 -527 -415 -521
rect -449 -595 -415 -593
rect -449 -631 -415 -629
rect -449 -703 -415 -697
rect -449 -775 -415 -765
rect -449 -847 -415 -833
rect -449 -919 -415 -901
rect -449 -991 -415 -969
rect -449 -1063 -415 -1037
rect -449 -1135 -415 -1105
rect -449 -1207 -415 -1173
rect -449 -1275 -415 -1241
rect -449 -1343 -415 -1313
rect -449 -1411 -415 -1385
rect -449 -1479 -415 -1457
rect -449 -1547 -415 -1529
rect -449 -1615 -415 -1601
rect -449 -1683 -415 -1673
rect -449 -1751 -415 -1745
rect -449 -1819 -415 -1817
rect -449 -1855 -415 -1853
rect -449 -1927 -415 -1921
rect -449 -1999 -415 -1989
rect -449 -2071 -415 -2057
rect -449 -2143 -415 -2125
rect -449 -2215 -415 -2193
rect -449 -2287 -415 -2261
rect -449 -2359 -415 -2329
rect -449 -2431 -415 -2397
rect -449 -2504 -415 -2465
rect -341 2465 -307 2504
rect -341 2397 -307 2431
rect -341 2329 -307 2359
rect -341 2261 -307 2287
rect -341 2193 -307 2215
rect -341 2125 -307 2143
rect -341 2057 -307 2071
rect -341 1989 -307 1999
rect -341 1921 -307 1927
rect -341 1853 -307 1855
rect -341 1817 -307 1819
rect -341 1745 -307 1751
rect -341 1673 -307 1683
rect -341 1601 -307 1615
rect -341 1529 -307 1547
rect -341 1457 -307 1479
rect -341 1385 -307 1411
rect -341 1313 -307 1343
rect -341 1241 -307 1275
rect -341 1173 -307 1207
rect -341 1105 -307 1135
rect -341 1037 -307 1063
rect -341 969 -307 991
rect -341 901 -307 919
rect -341 833 -307 847
rect -341 765 -307 775
rect -341 697 -307 703
rect -341 629 -307 631
rect -341 593 -307 595
rect -341 521 -307 527
rect -341 449 -307 459
rect -341 377 -307 391
rect -341 305 -307 323
rect -341 233 -307 255
rect -341 161 -307 187
rect -341 89 -307 119
rect -341 17 -307 51
rect -341 -51 -307 -17
rect -341 -119 -307 -89
rect -341 -187 -307 -161
rect -341 -255 -307 -233
rect -341 -323 -307 -305
rect -341 -391 -307 -377
rect -341 -459 -307 -449
rect -341 -527 -307 -521
rect -341 -595 -307 -593
rect -341 -631 -307 -629
rect -341 -703 -307 -697
rect -341 -775 -307 -765
rect -341 -847 -307 -833
rect -341 -919 -307 -901
rect -341 -991 -307 -969
rect -341 -1063 -307 -1037
rect -341 -1135 -307 -1105
rect -341 -1207 -307 -1173
rect -341 -1275 -307 -1241
rect -341 -1343 -307 -1313
rect -341 -1411 -307 -1385
rect -341 -1479 -307 -1457
rect -341 -1547 -307 -1529
rect -341 -1615 -307 -1601
rect -341 -1683 -307 -1673
rect -341 -1751 -307 -1745
rect -341 -1819 -307 -1817
rect -341 -1855 -307 -1853
rect -341 -1927 -307 -1921
rect -341 -1999 -307 -1989
rect -341 -2071 -307 -2057
rect -341 -2143 -307 -2125
rect -341 -2215 -307 -2193
rect -341 -2287 -307 -2261
rect -341 -2359 -307 -2329
rect -341 -2431 -307 -2397
rect -341 -2504 -307 -2465
rect -233 2465 -199 2504
rect -233 2397 -199 2431
rect -233 2329 -199 2359
rect -233 2261 -199 2287
rect -233 2193 -199 2215
rect -233 2125 -199 2143
rect -233 2057 -199 2071
rect -233 1989 -199 1999
rect -233 1921 -199 1927
rect -233 1853 -199 1855
rect -233 1817 -199 1819
rect -233 1745 -199 1751
rect -233 1673 -199 1683
rect -233 1601 -199 1615
rect -233 1529 -199 1547
rect -233 1457 -199 1479
rect -233 1385 -199 1411
rect -233 1313 -199 1343
rect -233 1241 -199 1275
rect -233 1173 -199 1207
rect -233 1105 -199 1135
rect -233 1037 -199 1063
rect -233 969 -199 991
rect -233 901 -199 919
rect -233 833 -199 847
rect -233 765 -199 775
rect -233 697 -199 703
rect -233 629 -199 631
rect -233 593 -199 595
rect -233 521 -199 527
rect -233 449 -199 459
rect -233 377 -199 391
rect -233 305 -199 323
rect -233 233 -199 255
rect -233 161 -199 187
rect -233 89 -199 119
rect -233 17 -199 51
rect -233 -51 -199 -17
rect -233 -119 -199 -89
rect -233 -187 -199 -161
rect -233 -255 -199 -233
rect -233 -323 -199 -305
rect -233 -391 -199 -377
rect -233 -459 -199 -449
rect -233 -527 -199 -521
rect -233 -595 -199 -593
rect -233 -631 -199 -629
rect -233 -703 -199 -697
rect -233 -775 -199 -765
rect -233 -847 -199 -833
rect -233 -919 -199 -901
rect -233 -991 -199 -969
rect -233 -1063 -199 -1037
rect -233 -1135 -199 -1105
rect -233 -1207 -199 -1173
rect -233 -1275 -199 -1241
rect -233 -1343 -199 -1313
rect -233 -1411 -199 -1385
rect -233 -1479 -199 -1457
rect -233 -1547 -199 -1529
rect -233 -1615 -199 -1601
rect -233 -1683 -199 -1673
rect -233 -1751 -199 -1745
rect -233 -1819 -199 -1817
rect -233 -1855 -199 -1853
rect -233 -1927 -199 -1921
rect -233 -1999 -199 -1989
rect -233 -2071 -199 -2057
rect -233 -2143 -199 -2125
rect -233 -2215 -199 -2193
rect -233 -2287 -199 -2261
rect -233 -2359 -199 -2329
rect -233 -2431 -199 -2397
rect -233 -2504 -199 -2465
rect -125 2465 -91 2504
rect -125 2397 -91 2431
rect -125 2329 -91 2359
rect -125 2261 -91 2287
rect -125 2193 -91 2215
rect -125 2125 -91 2143
rect -125 2057 -91 2071
rect -125 1989 -91 1999
rect -125 1921 -91 1927
rect -125 1853 -91 1855
rect -125 1817 -91 1819
rect -125 1745 -91 1751
rect -125 1673 -91 1683
rect -125 1601 -91 1615
rect -125 1529 -91 1547
rect -125 1457 -91 1479
rect -125 1385 -91 1411
rect -125 1313 -91 1343
rect -125 1241 -91 1275
rect -125 1173 -91 1207
rect -125 1105 -91 1135
rect -125 1037 -91 1063
rect -125 969 -91 991
rect -125 901 -91 919
rect -125 833 -91 847
rect -125 765 -91 775
rect -125 697 -91 703
rect -125 629 -91 631
rect -125 593 -91 595
rect -125 521 -91 527
rect -125 449 -91 459
rect -125 377 -91 391
rect -125 305 -91 323
rect -125 233 -91 255
rect -125 161 -91 187
rect -125 89 -91 119
rect -125 17 -91 51
rect -125 -51 -91 -17
rect -125 -119 -91 -89
rect -125 -187 -91 -161
rect -125 -255 -91 -233
rect -125 -323 -91 -305
rect -125 -391 -91 -377
rect -125 -459 -91 -449
rect -125 -527 -91 -521
rect -125 -595 -91 -593
rect -125 -631 -91 -629
rect -125 -703 -91 -697
rect -125 -775 -91 -765
rect -125 -847 -91 -833
rect -125 -919 -91 -901
rect -125 -991 -91 -969
rect -125 -1063 -91 -1037
rect -125 -1135 -91 -1105
rect -125 -1207 -91 -1173
rect -125 -1275 -91 -1241
rect -125 -1343 -91 -1313
rect -125 -1411 -91 -1385
rect -125 -1479 -91 -1457
rect -125 -1547 -91 -1529
rect -125 -1615 -91 -1601
rect -125 -1683 -91 -1673
rect -125 -1751 -91 -1745
rect -125 -1819 -91 -1817
rect -125 -1855 -91 -1853
rect -125 -1927 -91 -1921
rect -125 -1999 -91 -1989
rect -125 -2071 -91 -2057
rect -125 -2143 -91 -2125
rect -125 -2215 -91 -2193
rect -125 -2287 -91 -2261
rect -125 -2359 -91 -2329
rect -125 -2431 -91 -2397
rect -125 -2504 -91 -2465
rect -17 2465 17 2504
rect -17 2397 17 2431
rect -17 2329 17 2359
rect -17 2261 17 2287
rect -17 2193 17 2215
rect -17 2125 17 2143
rect -17 2057 17 2071
rect -17 1989 17 1999
rect -17 1921 17 1927
rect -17 1853 17 1855
rect -17 1817 17 1819
rect -17 1745 17 1751
rect -17 1673 17 1683
rect -17 1601 17 1615
rect -17 1529 17 1547
rect -17 1457 17 1479
rect -17 1385 17 1411
rect -17 1313 17 1343
rect -17 1241 17 1275
rect -17 1173 17 1207
rect -17 1105 17 1135
rect -17 1037 17 1063
rect -17 969 17 991
rect -17 901 17 919
rect -17 833 17 847
rect -17 765 17 775
rect -17 697 17 703
rect -17 629 17 631
rect -17 593 17 595
rect -17 521 17 527
rect -17 449 17 459
rect -17 377 17 391
rect -17 305 17 323
rect -17 233 17 255
rect -17 161 17 187
rect -17 89 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -89
rect -17 -187 17 -161
rect -17 -255 17 -233
rect -17 -323 17 -305
rect -17 -391 17 -377
rect -17 -459 17 -449
rect -17 -527 17 -521
rect -17 -595 17 -593
rect -17 -631 17 -629
rect -17 -703 17 -697
rect -17 -775 17 -765
rect -17 -847 17 -833
rect -17 -919 17 -901
rect -17 -991 17 -969
rect -17 -1063 17 -1037
rect -17 -1135 17 -1105
rect -17 -1207 17 -1173
rect -17 -1275 17 -1241
rect -17 -1343 17 -1313
rect -17 -1411 17 -1385
rect -17 -1479 17 -1457
rect -17 -1547 17 -1529
rect -17 -1615 17 -1601
rect -17 -1683 17 -1673
rect -17 -1751 17 -1745
rect -17 -1819 17 -1817
rect -17 -1855 17 -1853
rect -17 -1927 17 -1921
rect -17 -1999 17 -1989
rect -17 -2071 17 -2057
rect -17 -2143 17 -2125
rect -17 -2215 17 -2193
rect -17 -2287 17 -2261
rect -17 -2359 17 -2329
rect -17 -2431 17 -2397
rect -17 -2504 17 -2465
rect 91 2465 125 2504
rect 91 2397 125 2431
rect 91 2329 125 2359
rect 91 2261 125 2287
rect 91 2193 125 2215
rect 91 2125 125 2143
rect 91 2057 125 2071
rect 91 1989 125 1999
rect 91 1921 125 1927
rect 91 1853 125 1855
rect 91 1817 125 1819
rect 91 1745 125 1751
rect 91 1673 125 1683
rect 91 1601 125 1615
rect 91 1529 125 1547
rect 91 1457 125 1479
rect 91 1385 125 1411
rect 91 1313 125 1343
rect 91 1241 125 1275
rect 91 1173 125 1207
rect 91 1105 125 1135
rect 91 1037 125 1063
rect 91 969 125 991
rect 91 901 125 919
rect 91 833 125 847
rect 91 765 125 775
rect 91 697 125 703
rect 91 629 125 631
rect 91 593 125 595
rect 91 521 125 527
rect 91 449 125 459
rect 91 377 125 391
rect 91 305 125 323
rect 91 233 125 255
rect 91 161 125 187
rect 91 89 125 119
rect 91 17 125 51
rect 91 -51 125 -17
rect 91 -119 125 -89
rect 91 -187 125 -161
rect 91 -255 125 -233
rect 91 -323 125 -305
rect 91 -391 125 -377
rect 91 -459 125 -449
rect 91 -527 125 -521
rect 91 -595 125 -593
rect 91 -631 125 -629
rect 91 -703 125 -697
rect 91 -775 125 -765
rect 91 -847 125 -833
rect 91 -919 125 -901
rect 91 -991 125 -969
rect 91 -1063 125 -1037
rect 91 -1135 125 -1105
rect 91 -1207 125 -1173
rect 91 -1275 125 -1241
rect 91 -1343 125 -1313
rect 91 -1411 125 -1385
rect 91 -1479 125 -1457
rect 91 -1547 125 -1529
rect 91 -1615 125 -1601
rect 91 -1683 125 -1673
rect 91 -1751 125 -1745
rect 91 -1819 125 -1817
rect 91 -1855 125 -1853
rect 91 -1927 125 -1921
rect 91 -1999 125 -1989
rect 91 -2071 125 -2057
rect 91 -2143 125 -2125
rect 91 -2215 125 -2193
rect 91 -2287 125 -2261
rect 91 -2359 125 -2329
rect 91 -2431 125 -2397
rect 91 -2504 125 -2465
rect 199 2465 233 2504
rect 199 2397 233 2431
rect 199 2329 233 2359
rect 199 2261 233 2287
rect 199 2193 233 2215
rect 199 2125 233 2143
rect 199 2057 233 2071
rect 199 1989 233 1999
rect 199 1921 233 1927
rect 199 1853 233 1855
rect 199 1817 233 1819
rect 199 1745 233 1751
rect 199 1673 233 1683
rect 199 1601 233 1615
rect 199 1529 233 1547
rect 199 1457 233 1479
rect 199 1385 233 1411
rect 199 1313 233 1343
rect 199 1241 233 1275
rect 199 1173 233 1207
rect 199 1105 233 1135
rect 199 1037 233 1063
rect 199 969 233 991
rect 199 901 233 919
rect 199 833 233 847
rect 199 765 233 775
rect 199 697 233 703
rect 199 629 233 631
rect 199 593 233 595
rect 199 521 233 527
rect 199 449 233 459
rect 199 377 233 391
rect 199 305 233 323
rect 199 233 233 255
rect 199 161 233 187
rect 199 89 233 119
rect 199 17 233 51
rect 199 -51 233 -17
rect 199 -119 233 -89
rect 199 -187 233 -161
rect 199 -255 233 -233
rect 199 -323 233 -305
rect 199 -391 233 -377
rect 199 -459 233 -449
rect 199 -527 233 -521
rect 199 -595 233 -593
rect 199 -631 233 -629
rect 199 -703 233 -697
rect 199 -775 233 -765
rect 199 -847 233 -833
rect 199 -919 233 -901
rect 199 -991 233 -969
rect 199 -1063 233 -1037
rect 199 -1135 233 -1105
rect 199 -1207 233 -1173
rect 199 -1275 233 -1241
rect 199 -1343 233 -1313
rect 199 -1411 233 -1385
rect 199 -1479 233 -1457
rect 199 -1547 233 -1529
rect 199 -1615 233 -1601
rect 199 -1683 233 -1673
rect 199 -1751 233 -1745
rect 199 -1819 233 -1817
rect 199 -1855 233 -1853
rect 199 -1927 233 -1921
rect 199 -1999 233 -1989
rect 199 -2071 233 -2057
rect 199 -2143 233 -2125
rect 199 -2215 233 -2193
rect 199 -2287 233 -2261
rect 199 -2359 233 -2329
rect 199 -2431 233 -2397
rect 199 -2504 233 -2465
rect 307 2465 341 2504
rect 307 2397 341 2431
rect 307 2329 341 2359
rect 307 2261 341 2287
rect 307 2193 341 2215
rect 307 2125 341 2143
rect 307 2057 341 2071
rect 307 1989 341 1999
rect 307 1921 341 1927
rect 307 1853 341 1855
rect 307 1817 341 1819
rect 307 1745 341 1751
rect 307 1673 341 1683
rect 307 1601 341 1615
rect 307 1529 341 1547
rect 307 1457 341 1479
rect 307 1385 341 1411
rect 307 1313 341 1343
rect 307 1241 341 1275
rect 307 1173 341 1207
rect 307 1105 341 1135
rect 307 1037 341 1063
rect 307 969 341 991
rect 307 901 341 919
rect 307 833 341 847
rect 307 765 341 775
rect 307 697 341 703
rect 307 629 341 631
rect 307 593 341 595
rect 307 521 341 527
rect 307 449 341 459
rect 307 377 341 391
rect 307 305 341 323
rect 307 233 341 255
rect 307 161 341 187
rect 307 89 341 119
rect 307 17 341 51
rect 307 -51 341 -17
rect 307 -119 341 -89
rect 307 -187 341 -161
rect 307 -255 341 -233
rect 307 -323 341 -305
rect 307 -391 341 -377
rect 307 -459 341 -449
rect 307 -527 341 -521
rect 307 -595 341 -593
rect 307 -631 341 -629
rect 307 -703 341 -697
rect 307 -775 341 -765
rect 307 -847 341 -833
rect 307 -919 341 -901
rect 307 -991 341 -969
rect 307 -1063 341 -1037
rect 307 -1135 341 -1105
rect 307 -1207 341 -1173
rect 307 -1275 341 -1241
rect 307 -1343 341 -1313
rect 307 -1411 341 -1385
rect 307 -1479 341 -1457
rect 307 -1547 341 -1529
rect 307 -1615 341 -1601
rect 307 -1683 341 -1673
rect 307 -1751 341 -1745
rect 307 -1819 341 -1817
rect 307 -1855 341 -1853
rect 307 -1927 341 -1921
rect 307 -1999 341 -1989
rect 307 -2071 341 -2057
rect 307 -2143 341 -2125
rect 307 -2215 341 -2193
rect 307 -2287 341 -2261
rect 307 -2359 341 -2329
rect 307 -2431 341 -2397
rect 307 -2504 341 -2465
rect 415 2465 449 2504
rect 415 2397 449 2431
rect 415 2329 449 2359
rect 415 2261 449 2287
rect 415 2193 449 2215
rect 415 2125 449 2143
rect 415 2057 449 2071
rect 415 1989 449 1999
rect 415 1921 449 1927
rect 415 1853 449 1855
rect 415 1817 449 1819
rect 415 1745 449 1751
rect 415 1673 449 1683
rect 415 1601 449 1615
rect 415 1529 449 1547
rect 415 1457 449 1479
rect 415 1385 449 1411
rect 415 1313 449 1343
rect 415 1241 449 1275
rect 415 1173 449 1207
rect 415 1105 449 1135
rect 415 1037 449 1063
rect 415 969 449 991
rect 415 901 449 919
rect 415 833 449 847
rect 415 765 449 775
rect 415 697 449 703
rect 415 629 449 631
rect 415 593 449 595
rect 415 521 449 527
rect 415 449 449 459
rect 415 377 449 391
rect 415 305 449 323
rect 415 233 449 255
rect 415 161 449 187
rect 415 89 449 119
rect 415 17 449 51
rect 415 -51 449 -17
rect 415 -119 449 -89
rect 415 -187 449 -161
rect 415 -255 449 -233
rect 415 -323 449 -305
rect 415 -391 449 -377
rect 415 -459 449 -449
rect 415 -527 449 -521
rect 415 -595 449 -593
rect 415 -631 449 -629
rect 415 -703 449 -697
rect 415 -775 449 -765
rect 415 -847 449 -833
rect 415 -919 449 -901
rect 415 -991 449 -969
rect 415 -1063 449 -1037
rect 415 -1135 449 -1105
rect 415 -1207 449 -1173
rect 415 -1275 449 -1241
rect 415 -1343 449 -1313
rect 415 -1411 449 -1385
rect 415 -1479 449 -1457
rect 415 -1547 449 -1529
rect 415 -1615 449 -1601
rect 415 -1683 449 -1673
rect 415 -1751 449 -1745
rect 415 -1819 449 -1817
rect 415 -1855 449 -1853
rect 415 -1927 449 -1921
rect 415 -1999 449 -1989
rect 415 -2071 449 -2057
rect 415 -2143 449 -2125
rect 415 -2215 449 -2193
rect 415 -2287 449 -2261
rect 415 -2359 449 -2329
rect 415 -2431 449 -2397
rect 415 -2504 449 -2465
rect 529 2499 563 2533
rect 529 2431 563 2465
rect 529 2363 563 2397
rect 529 2295 563 2329
rect 529 2227 563 2261
rect 529 2159 563 2193
rect 529 2091 563 2125
rect 529 2023 563 2057
rect 529 1955 563 1989
rect 529 1887 563 1921
rect 529 1819 563 1853
rect 529 1751 563 1785
rect 529 1683 563 1717
rect 529 1615 563 1649
rect 529 1547 563 1581
rect 529 1479 563 1513
rect 529 1411 563 1445
rect 529 1343 563 1377
rect 529 1275 563 1309
rect 529 1207 563 1241
rect 529 1139 563 1173
rect 529 1071 563 1105
rect 529 1003 563 1037
rect 529 935 563 969
rect 529 867 563 901
rect 529 799 563 833
rect 529 731 563 765
rect 529 663 563 697
rect 529 595 563 629
rect 529 527 563 561
rect 529 459 563 493
rect 529 391 563 425
rect 529 323 563 357
rect 529 255 563 289
rect 529 187 563 221
rect 529 119 563 153
rect 529 51 563 85
rect 529 -17 563 17
rect 529 -85 563 -51
rect 529 -153 563 -119
rect 529 -221 563 -187
rect 529 -289 563 -255
rect 529 -357 563 -323
rect 529 -425 563 -391
rect 529 -493 563 -459
rect 529 -561 563 -527
rect 529 -629 563 -595
rect 529 -697 563 -663
rect 529 -765 563 -731
rect 529 -833 563 -799
rect 529 -901 563 -867
rect 529 -969 563 -935
rect 529 -1037 563 -1003
rect 529 -1105 563 -1071
rect 529 -1173 563 -1139
rect 529 -1241 563 -1207
rect 529 -1309 563 -1275
rect 529 -1377 563 -1343
rect 529 -1445 563 -1411
rect 529 -1513 563 -1479
rect 529 -1581 563 -1547
rect 529 -1649 563 -1615
rect 529 -1717 563 -1683
rect 529 -1785 563 -1751
rect 529 -1853 563 -1819
rect 529 -1921 563 -1887
rect 529 -1989 563 -1955
rect 529 -2057 563 -2023
rect 529 -2125 563 -2091
rect 529 -2193 563 -2159
rect 529 -2261 563 -2227
rect 529 -2329 563 -2295
rect 529 -2397 563 -2363
rect 529 -2465 563 -2431
rect 529 -2533 563 -2499
rect -563 -2649 -529 -2567
rect -411 -2581 -395 -2547
rect -361 -2581 -345 -2547
rect -195 -2581 -179 -2547
rect -145 -2581 -129 -2547
rect 21 -2581 37 -2547
rect 71 -2581 87 -2547
rect 237 -2581 253 -2547
rect 287 -2581 303 -2547
rect 529 -2649 563 -2567
rect -563 -2683 -459 -2649
rect -425 -2683 -391 -2649
rect -357 -2683 -323 -2649
rect -289 -2683 -255 -2649
rect -221 -2683 -187 -2649
rect -153 -2683 -119 -2649
rect -85 -2683 -51 -2649
rect -17 -2683 17 -2649
rect 51 -2683 85 -2649
rect 119 -2683 153 -2649
rect 187 -2683 221 -2649
rect 255 -2683 289 -2649
rect 323 -2683 357 -2649
rect 391 -2683 425 -2649
rect 459 -2683 563 -2649
<< viali >>
rect -287 2547 -253 2581
rect -71 2547 -37 2581
rect 145 2547 179 2581
rect 361 2547 395 2581
rect -449 2431 -415 2465
rect -449 2363 -415 2393
rect -449 2359 -415 2363
rect -449 2295 -415 2321
rect -449 2287 -415 2295
rect -449 2227 -415 2249
rect -449 2215 -415 2227
rect -449 2159 -415 2177
rect -449 2143 -415 2159
rect -449 2091 -415 2105
rect -449 2071 -415 2091
rect -449 2023 -415 2033
rect -449 1999 -415 2023
rect -449 1955 -415 1961
rect -449 1927 -415 1955
rect -449 1887 -415 1889
rect -449 1855 -415 1887
rect -449 1785 -415 1817
rect -449 1783 -415 1785
rect -449 1717 -415 1745
rect -449 1711 -415 1717
rect -449 1649 -415 1673
rect -449 1639 -415 1649
rect -449 1581 -415 1601
rect -449 1567 -415 1581
rect -449 1513 -415 1529
rect -449 1495 -415 1513
rect -449 1445 -415 1457
rect -449 1423 -415 1445
rect -449 1377 -415 1385
rect -449 1351 -415 1377
rect -449 1309 -415 1313
rect -449 1279 -415 1309
rect -449 1207 -415 1241
rect -449 1139 -415 1169
rect -449 1135 -415 1139
rect -449 1071 -415 1097
rect -449 1063 -415 1071
rect -449 1003 -415 1025
rect -449 991 -415 1003
rect -449 935 -415 953
rect -449 919 -415 935
rect -449 867 -415 881
rect -449 847 -415 867
rect -449 799 -415 809
rect -449 775 -415 799
rect -449 731 -415 737
rect -449 703 -415 731
rect -449 663 -415 665
rect -449 631 -415 663
rect -449 561 -415 593
rect -449 559 -415 561
rect -449 493 -415 521
rect -449 487 -415 493
rect -449 425 -415 449
rect -449 415 -415 425
rect -449 357 -415 377
rect -449 343 -415 357
rect -449 289 -415 305
rect -449 271 -415 289
rect -449 221 -415 233
rect -449 199 -415 221
rect -449 153 -415 161
rect -449 127 -415 153
rect -449 85 -415 89
rect -449 55 -415 85
rect -449 -17 -415 17
rect -449 -85 -415 -55
rect -449 -89 -415 -85
rect -449 -153 -415 -127
rect -449 -161 -415 -153
rect -449 -221 -415 -199
rect -449 -233 -415 -221
rect -449 -289 -415 -271
rect -449 -305 -415 -289
rect -449 -357 -415 -343
rect -449 -377 -415 -357
rect -449 -425 -415 -415
rect -449 -449 -415 -425
rect -449 -493 -415 -487
rect -449 -521 -415 -493
rect -449 -561 -415 -559
rect -449 -593 -415 -561
rect -449 -663 -415 -631
rect -449 -665 -415 -663
rect -449 -731 -415 -703
rect -449 -737 -415 -731
rect -449 -799 -415 -775
rect -449 -809 -415 -799
rect -449 -867 -415 -847
rect -449 -881 -415 -867
rect -449 -935 -415 -919
rect -449 -953 -415 -935
rect -449 -1003 -415 -991
rect -449 -1025 -415 -1003
rect -449 -1071 -415 -1063
rect -449 -1097 -415 -1071
rect -449 -1139 -415 -1135
rect -449 -1169 -415 -1139
rect -449 -1241 -415 -1207
rect -449 -1309 -415 -1279
rect -449 -1313 -415 -1309
rect -449 -1377 -415 -1351
rect -449 -1385 -415 -1377
rect -449 -1445 -415 -1423
rect -449 -1457 -415 -1445
rect -449 -1513 -415 -1495
rect -449 -1529 -415 -1513
rect -449 -1581 -415 -1567
rect -449 -1601 -415 -1581
rect -449 -1649 -415 -1639
rect -449 -1673 -415 -1649
rect -449 -1717 -415 -1711
rect -449 -1745 -415 -1717
rect -449 -1785 -415 -1783
rect -449 -1817 -415 -1785
rect -449 -1887 -415 -1855
rect -449 -1889 -415 -1887
rect -449 -1955 -415 -1927
rect -449 -1961 -415 -1955
rect -449 -2023 -415 -1999
rect -449 -2033 -415 -2023
rect -449 -2091 -415 -2071
rect -449 -2105 -415 -2091
rect -449 -2159 -415 -2143
rect -449 -2177 -415 -2159
rect -449 -2227 -415 -2215
rect -449 -2249 -415 -2227
rect -449 -2295 -415 -2287
rect -449 -2321 -415 -2295
rect -449 -2363 -415 -2359
rect -449 -2393 -415 -2363
rect -449 -2465 -415 -2431
rect -341 2431 -307 2465
rect -341 2363 -307 2393
rect -341 2359 -307 2363
rect -341 2295 -307 2321
rect -341 2287 -307 2295
rect -341 2227 -307 2249
rect -341 2215 -307 2227
rect -341 2159 -307 2177
rect -341 2143 -307 2159
rect -341 2091 -307 2105
rect -341 2071 -307 2091
rect -341 2023 -307 2033
rect -341 1999 -307 2023
rect -341 1955 -307 1961
rect -341 1927 -307 1955
rect -341 1887 -307 1889
rect -341 1855 -307 1887
rect -341 1785 -307 1817
rect -341 1783 -307 1785
rect -341 1717 -307 1745
rect -341 1711 -307 1717
rect -341 1649 -307 1673
rect -341 1639 -307 1649
rect -341 1581 -307 1601
rect -341 1567 -307 1581
rect -341 1513 -307 1529
rect -341 1495 -307 1513
rect -341 1445 -307 1457
rect -341 1423 -307 1445
rect -341 1377 -307 1385
rect -341 1351 -307 1377
rect -341 1309 -307 1313
rect -341 1279 -307 1309
rect -341 1207 -307 1241
rect -341 1139 -307 1169
rect -341 1135 -307 1139
rect -341 1071 -307 1097
rect -341 1063 -307 1071
rect -341 1003 -307 1025
rect -341 991 -307 1003
rect -341 935 -307 953
rect -341 919 -307 935
rect -341 867 -307 881
rect -341 847 -307 867
rect -341 799 -307 809
rect -341 775 -307 799
rect -341 731 -307 737
rect -341 703 -307 731
rect -341 663 -307 665
rect -341 631 -307 663
rect -341 561 -307 593
rect -341 559 -307 561
rect -341 493 -307 521
rect -341 487 -307 493
rect -341 425 -307 449
rect -341 415 -307 425
rect -341 357 -307 377
rect -341 343 -307 357
rect -341 289 -307 305
rect -341 271 -307 289
rect -341 221 -307 233
rect -341 199 -307 221
rect -341 153 -307 161
rect -341 127 -307 153
rect -341 85 -307 89
rect -341 55 -307 85
rect -341 -17 -307 17
rect -341 -85 -307 -55
rect -341 -89 -307 -85
rect -341 -153 -307 -127
rect -341 -161 -307 -153
rect -341 -221 -307 -199
rect -341 -233 -307 -221
rect -341 -289 -307 -271
rect -341 -305 -307 -289
rect -341 -357 -307 -343
rect -341 -377 -307 -357
rect -341 -425 -307 -415
rect -341 -449 -307 -425
rect -341 -493 -307 -487
rect -341 -521 -307 -493
rect -341 -561 -307 -559
rect -341 -593 -307 -561
rect -341 -663 -307 -631
rect -341 -665 -307 -663
rect -341 -731 -307 -703
rect -341 -737 -307 -731
rect -341 -799 -307 -775
rect -341 -809 -307 -799
rect -341 -867 -307 -847
rect -341 -881 -307 -867
rect -341 -935 -307 -919
rect -341 -953 -307 -935
rect -341 -1003 -307 -991
rect -341 -1025 -307 -1003
rect -341 -1071 -307 -1063
rect -341 -1097 -307 -1071
rect -341 -1139 -307 -1135
rect -341 -1169 -307 -1139
rect -341 -1241 -307 -1207
rect -341 -1309 -307 -1279
rect -341 -1313 -307 -1309
rect -341 -1377 -307 -1351
rect -341 -1385 -307 -1377
rect -341 -1445 -307 -1423
rect -341 -1457 -307 -1445
rect -341 -1513 -307 -1495
rect -341 -1529 -307 -1513
rect -341 -1581 -307 -1567
rect -341 -1601 -307 -1581
rect -341 -1649 -307 -1639
rect -341 -1673 -307 -1649
rect -341 -1717 -307 -1711
rect -341 -1745 -307 -1717
rect -341 -1785 -307 -1783
rect -341 -1817 -307 -1785
rect -341 -1887 -307 -1855
rect -341 -1889 -307 -1887
rect -341 -1955 -307 -1927
rect -341 -1961 -307 -1955
rect -341 -2023 -307 -1999
rect -341 -2033 -307 -2023
rect -341 -2091 -307 -2071
rect -341 -2105 -307 -2091
rect -341 -2159 -307 -2143
rect -341 -2177 -307 -2159
rect -341 -2227 -307 -2215
rect -341 -2249 -307 -2227
rect -341 -2295 -307 -2287
rect -341 -2321 -307 -2295
rect -341 -2363 -307 -2359
rect -341 -2393 -307 -2363
rect -341 -2465 -307 -2431
rect -233 2431 -199 2465
rect -233 2363 -199 2393
rect -233 2359 -199 2363
rect -233 2295 -199 2321
rect -233 2287 -199 2295
rect -233 2227 -199 2249
rect -233 2215 -199 2227
rect -233 2159 -199 2177
rect -233 2143 -199 2159
rect -233 2091 -199 2105
rect -233 2071 -199 2091
rect -233 2023 -199 2033
rect -233 1999 -199 2023
rect -233 1955 -199 1961
rect -233 1927 -199 1955
rect -233 1887 -199 1889
rect -233 1855 -199 1887
rect -233 1785 -199 1817
rect -233 1783 -199 1785
rect -233 1717 -199 1745
rect -233 1711 -199 1717
rect -233 1649 -199 1673
rect -233 1639 -199 1649
rect -233 1581 -199 1601
rect -233 1567 -199 1581
rect -233 1513 -199 1529
rect -233 1495 -199 1513
rect -233 1445 -199 1457
rect -233 1423 -199 1445
rect -233 1377 -199 1385
rect -233 1351 -199 1377
rect -233 1309 -199 1313
rect -233 1279 -199 1309
rect -233 1207 -199 1241
rect -233 1139 -199 1169
rect -233 1135 -199 1139
rect -233 1071 -199 1097
rect -233 1063 -199 1071
rect -233 1003 -199 1025
rect -233 991 -199 1003
rect -233 935 -199 953
rect -233 919 -199 935
rect -233 867 -199 881
rect -233 847 -199 867
rect -233 799 -199 809
rect -233 775 -199 799
rect -233 731 -199 737
rect -233 703 -199 731
rect -233 663 -199 665
rect -233 631 -199 663
rect -233 561 -199 593
rect -233 559 -199 561
rect -233 493 -199 521
rect -233 487 -199 493
rect -233 425 -199 449
rect -233 415 -199 425
rect -233 357 -199 377
rect -233 343 -199 357
rect -233 289 -199 305
rect -233 271 -199 289
rect -233 221 -199 233
rect -233 199 -199 221
rect -233 153 -199 161
rect -233 127 -199 153
rect -233 85 -199 89
rect -233 55 -199 85
rect -233 -17 -199 17
rect -233 -85 -199 -55
rect -233 -89 -199 -85
rect -233 -153 -199 -127
rect -233 -161 -199 -153
rect -233 -221 -199 -199
rect -233 -233 -199 -221
rect -233 -289 -199 -271
rect -233 -305 -199 -289
rect -233 -357 -199 -343
rect -233 -377 -199 -357
rect -233 -425 -199 -415
rect -233 -449 -199 -425
rect -233 -493 -199 -487
rect -233 -521 -199 -493
rect -233 -561 -199 -559
rect -233 -593 -199 -561
rect -233 -663 -199 -631
rect -233 -665 -199 -663
rect -233 -731 -199 -703
rect -233 -737 -199 -731
rect -233 -799 -199 -775
rect -233 -809 -199 -799
rect -233 -867 -199 -847
rect -233 -881 -199 -867
rect -233 -935 -199 -919
rect -233 -953 -199 -935
rect -233 -1003 -199 -991
rect -233 -1025 -199 -1003
rect -233 -1071 -199 -1063
rect -233 -1097 -199 -1071
rect -233 -1139 -199 -1135
rect -233 -1169 -199 -1139
rect -233 -1241 -199 -1207
rect -233 -1309 -199 -1279
rect -233 -1313 -199 -1309
rect -233 -1377 -199 -1351
rect -233 -1385 -199 -1377
rect -233 -1445 -199 -1423
rect -233 -1457 -199 -1445
rect -233 -1513 -199 -1495
rect -233 -1529 -199 -1513
rect -233 -1581 -199 -1567
rect -233 -1601 -199 -1581
rect -233 -1649 -199 -1639
rect -233 -1673 -199 -1649
rect -233 -1717 -199 -1711
rect -233 -1745 -199 -1717
rect -233 -1785 -199 -1783
rect -233 -1817 -199 -1785
rect -233 -1887 -199 -1855
rect -233 -1889 -199 -1887
rect -233 -1955 -199 -1927
rect -233 -1961 -199 -1955
rect -233 -2023 -199 -1999
rect -233 -2033 -199 -2023
rect -233 -2091 -199 -2071
rect -233 -2105 -199 -2091
rect -233 -2159 -199 -2143
rect -233 -2177 -199 -2159
rect -233 -2227 -199 -2215
rect -233 -2249 -199 -2227
rect -233 -2295 -199 -2287
rect -233 -2321 -199 -2295
rect -233 -2363 -199 -2359
rect -233 -2393 -199 -2363
rect -233 -2465 -199 -2431
rect -125 2431 -91 2465
rect -125 2363 -91 2393
rect -125 2359 -91 2363
rect -125 2295 -91 2321
rect -125 2287 -91 2295
rect -125 2227 -91 2249
rect -125 2215 -91 2227
rect -125 2159 -91 2177
rect -125 2143 -91 2159
rect -125 2091 -91 2105
rect -125 2071 -91 2091
rect -125 2023 -91 2033
rect -125 1999 -91 2023
rect -125 1955 -91 1961
rect -125 1927 -91 1955
rect -125 1887 -91 1889
rect -125 1855 -91 1887
rect -125 1785 -91 1817
rect -125 1783 -91 1785
rect -125 1717 -91 1745
rect -125 1711 -91 1717
rect -125 1649 -91 1673
rect -125 1639 -91 1649
rect -125 1581 -91 1601
rect -125 1567 -91 1581
rect -125 1513 -91 1529
rect -125 1495 -91 1513
rect -125 1445 -91 1457
rect -125 1423 -91 1445
rect -125 1377 -91 1385
rect -125 1351 -91 1377
rect -125 1309 -91 1313
rect -125 1279 -91 1309
rect -125 1207 -91 1241
rect -125 1139 -91 1169
rect -125 1135 -91 1139
rect -125 1071 -91 1097
rect -125 1063 -91 1071
rect -125 1003 -91 1025
rect -125 991 -91 1003
rect -125 935 -91 953
rect -125 919 -91 935
rect -125 867 -91 881
rect -125 847 -91 867
rect -125 799 -91 809
rect -125 775 -91 799
rect -125 731 -91 737
rect -125 703 -91 731
rect -125 663 -91 665
rect -125 631 -91 663
rect -125 561 -91 593
rect -125 559 -91 561
rect -125 493 -91 521
rect -125 487 -91 493
rect -125 425 -91 449
rect -125 415 -91 425
rect -125 357 -91 377
rect -125 343 -91 357
rect -125 289 -91 305
rect -125 271 -91 289
rect -125 221 -91 233
rect -125 199 -91 221
rect -125 153 -91 161
rect -125 127 -91 153
rect -125 85 -91 89
rect -125 55 -91 85
rect -125 -17 -91 17
rect -125 -85 -91 -55
rect -125 -89 -91 -85
rect -125 -153 -91 -127
rect -125 -161 -91 -153
rect -125 -221 -91 -199
rect -125 -233 -91 -221
rect -125 -289 -91 -271
rect -125 -305 -91 -289
rect -125 -357 -91 -343
rect -125 -377 -91 -357
rect -125 -425 -91 -415
rect -125 -449 -91 -425
rect -125 -493 -91 -487
rect -125 -521 -91 -493
rect -125 -561 -91 -559
rect -125 -593 -91 -561
rect -125 -663 -91 -631
rect -125 -665 -91 -663
rect -125 -731 -91 -703
rect -125 -737 -91 -731
rect -125 -799 -91 -775
rect -125 -809 -91 -799
rect -125 -867 -91 -847
rect -125 -881 -91 -867
rect -125 -935 -91 -919
rect -125 -953 -91 -935
rect -125 -1003 -91 -991
rect -125 -1025 -91 -1003
rect -125 -1071 -91 -1063
rect -125 -1097 -91 -1071
rect -125 -1139 -91 -1135
rect -125 -1169 -91 -1139
rect -125 -1241 -91 -1207
rect -125 -1309 -91 -1279
rect -125 -1313 -91 -1309
rect -125 -1377 -91 -1351
rect -125 -1385 -91 -1377
rect -125 -1445 -91 -1423
rect -125 -1457 -91 -1445
rect -125 -1513 -91 -1495
rect -125 -1529 -91 -1513
rect -125 -1581 -91 -1567
rect -125 -1601 -91 -1581
rect -125 -1649 -91 -1639
rect -125 -1673 -91 -1649
rect -125 -1717 -91 -1711
rect -125 -1745 -91 -1717
rect -125 -1785 -91 -1783
rect -125 -1817 -91 -1785
rect -125 -1887 -91 -1855
rect -125 -1889 -91 -1887
rect -125 -1955 -91 -1927
rect -125 -1961 -91 -1955
rect -125 -2023 -91 -1999
rect -125 -2033 -91 -2023
rect -125 -2091 -91 -2071
rect -125 -2105 -91 -2091
rect -125 -2159 -91 -2143
rect -125 -2177 -91 -2159
rect -125 -2227 -91 -2215
rect -125 -2249 -91 -2227
rect -125 -2295 -91 -2287
rect -125 -2321 -91 -2295
rect -125 -2363 -91 -2359
rect -125 -2393 -91 -2363
rect -125 -2465 -91 -2431
rect -17 2431 17 2465
rect -17 2363 17 2393
rect -17 2359 17 2363
rect -17 2295 17 2321
rect -17 2287 17 2295
rect -17 2227 17 2249
rect -17 2215 17 2227
rect -17 2159 17 2177
rect -17 2143 17 2159
rect -17 2091 17 2105
rect -17 2071 17 2091
rect -17 2023 17 2033
rect -17 1999 17 2023
rect -17 1955 17 1961
rect -17 1927 17 1955
rect -17 1887 17 1889
rect -17 1855 17 1887
rect -17 1785 17 1817
rect -17 1783 17 1785
rect -17 1717 17 1745
rect -17 1711 17 1717
rect -17 1649 17 1673
rect -17 1639 17 1649
rect -17 1581 17 1601
rect -17 1567 17 1581
rect -17 1513 17 1529
rect -17 1495 17 1513
rect -17 1445 17 1457
rect -17 1423 17 1445
rect -17 1377 17 1385
rect -17 1351 17 1377
rect -17 1309 17 1313
rect -17 1279 17 1309
rect -17 1207 17 1241
rect -17 1139 17 1169
rect -17 1135 17 1139
rect -17 1071 17 1097
rect -17 1063 17 1071
rect -17 1003 17 1025
rect -17 991 17 1003
rect -17 935 17 953
rect -17 919 17 935
rect -17 867 17 881
rect -17 847 17 867
rect -17 799 17 809
rect -17 775 17 799
rect -17 731 17 737
rect -17 703 17 731
rect -17 663 17 665
rect -17 631 17 663
rect -17 561 17 593
rect -17 559 17 561
rect -17 493 17 521
rect -17 487 17 493
rect -17 425 17 449
rect -17 415 17 425
rect -17 357 17 377
rect -17 343 17 357
rect -17 289 17 305
rect -17 271 17 289
rect -17 221 17 233
rect -17 199 17 221
rect -17 153 17 161
rect -17 127 17 153
rect -17 85 17 89
rect -17 55 17 85
rect -17 -17 17 17
rect -17 -85 17 -55
rect -17 -89 17 -85
rect -17 -153 17 -127
rect -17 -161 17 -153
rect -17 -221 17 -199
rect -17 -233 17 -221
rect -17 -289 17 -271
rect -17 -305 17 -289
rect -17 -357 17 -343
rect -17 -377 17 -357
rect -17 -425 17 -415
rect -17 -449 17 -425
rect -17 -493 17 -487
rect -17 -521 17 -493
rect -17 -561 17 -559
rect -17 -593 17 -561
rect -17 -663 17 -631
rect -17 -665 17 -663
rect -17 -731 17 -703
rect -17 -737 17 -731
rect -17 -799 17 -775
rect -17 -809 17 -799
rect -17 -867 17 -847
rect -17 -881 17 -867
rect -17 -935 17 -919
rect -17 -953 17 -935
rect -17 -1003 17 -991
rect -17 -1025 17 -1003
rect -17 -1071 17 -1063
rect -17 -1097 17 -1071
rect -17 -1139 17 -1135
rect -17 -1169 17 -1139
rect -17 -1241 17 -1207
rect -17 -1309 17 -1279
rect -17 -1313 17 -1309
rect -17 -1377 17 -1351
rect -17 -1385 17 -1377
rect -17 -1445 17 -1423
rect -17 -1457 17 -1445
rect -17 -1513 17 -1495
rect -17 -1529 17 -1513
rect -17 -1581 17 -1567
rect -17 -1601 17 -1581
rect -17 -1649 17 -1639
rect -17 -1673 17 -1649
rect -17 -1717 17 -1711
rect -17 -1745 17 -1717
rect -17 -1785 17 -1783
rect -17 -1817 17 -1785
rect -17 -1887 17 -1855
rect -17 -1889 17 -1887
rect -17 -1955 17 -1927
rect -17 -1961 17 -1955
rect -17 -2023 17 -1999
rect -17 -2033 17 -2023
rect -17 -2091 17 -2071
rect -17 -2105 17 -2091
rect -17 -2159 17 -2143
rect -17 -2177 17 -2159
rect -17 -2227 17 -2215
rect -17 -2249 17 -2227
rect -17 -2295 17 -2287
rect -17 -2321 17 -2295
rect -17 -2363 17 -2359
rect -17 -2393 17 -2363
rect -17 -2465 17 -2431
rect 91 2431 125 2465
rect 91 2363 125 2393
rect 91 2359 125 2363
rect 91 2295 125 2321
rect 91 2287 125 2295
rect 91 2227 125 2249
rect 91 2215 125 2227
rect 91 2159 125 2177
rect 91 2143 125 2159
rect 91 2091 125 2105
rect 91 2071 125 2091
rect 91 2023 125 2033
rect 91 1999 125 2023
rect 91 1955 125 1961
rect 91 1927 125 1955
rect 91 1887 125 1889
rect 91 1855 125 1887
rect 91 1785 125 1817
rect 91 1783 125 1785
rect 91 1717 125 1745
rect 91 1711 125 1717
rect 91 1649 125 1673
rect 91 1639 125 1649
rect 91 1581 125 1601
rect 91 1567 125 1581
rect 91 1513 125 1529
rect 91 1495 125 1513
rect 91 1445 125 1457
rect 91 1423 125 1445
rect 91 1377 125 1385
rect 91 1351 125 1377
rect 91 1309 125 1313
rect 91 1279 125 1309
rect 91 1207 125 1241
rect 91 1139 125 1169
rect 91 1135 125 1139
rect 91 1071 125 1097
rect 91 1063 125 1071
rect 91 1003 125 1025
rect 91 991 125 1003
rect 91 935 125 953
rect 91 919 125 935
rect 91 867 125 881
rect 91 847 125 867
rect 91 799 125 809
rect 91 775 125 799
rect 91 731 125 737
rect 91 703 125 731
rect 91 663 125 665
rect 91 631 125 663
rect 91 561 125 593
rect 91 559 125 561
rect 91 493 125 521
rect 91 487 125 493
rect 91 425 125 449
rect 91 415 125 425
rect 91 357 125 377
rect 91 343 125 357
rect 91 289 125 305
rect 91 271 125 289
rect 91 221 125 233
rect 91 199 125 221
rect 91 153 125 161
rect 91 127 125 153
rect 91 85 125 89
rect 91 55 125 85
rect 91 -17 125 17
rect 91 -85 125 -55
rect 91 -89 125 -85
rect 91 -153 125 -127
rect 91 -161 125 -153
rect 91 -221 125 -199
rect 91 -233 125 -221
rect 91 -289 125 -271
rect 91 -305 125 -289
rect 91 -357 125 -343
rect 91 -377 125 -357
rect 91 -425 125 -415
rect 91 -449 125 -425
rect 91 -493 125 -487
rect 91 -521 125 -493
rect 91 -561 125 -559
rect 91 -593 125 -561
rect 91 -663 125 -631
rect 91 -665 125 -663
rect 91 -731 125 -703
rect 91 -737 125 -731
rect 91 -799 125 -775
rect 91 -809 125 -799
rect 91 -867 125 -847
rect 91 -881 125 -867
rect 91 -935 125 -919
rect 91 -953 125 -935
rect 91 -1003 125 -991
rect 91 -1025 125 -1003
rect 91 -1071 125 -1063
rect 91 -1097 125 -1071
rect 91 -1139 125 -1135
rect 91 -1169 125 -1139
rect 91 -1241 125 -1207
rect 91 -1309 125 -1279
rect 91 -1313 125 -1309
rect 91 -1377 125 -1351
rect 91 -1385 125 -1377
rect 91 -1445 125 -1423
rect 91 -1457 125 -1445
rect 91 -1513 125 -1495
rect 91 -1529 125 -1513
rect 91 -1581 125 -1567
rect 91 -1601 125 -1581
rect 91 -1649 125 -1639
rect 91 -1673 125 -1649
rect 91 -1717 125 -1711
rect 91 -1745 125 -1717
rect 91 -1785 125 -1783
rect 91 -1817 125 -1785
rect 91 -1887 125 -1855
rect 91 -1889 125 -1887
rect 91 -1955 125 -1927
rect 91 -1961 125 -1955
rect 91 -2023 125 -1999
rect 91 -2033 125 -2023
rect 91 -2091 125 -2071
rect 91 -2105 125 -2091
rect 91 -2159 125 -2143
rect 91 -2177 125 -2159
rect 91 -2227 125 -2215
rect 91 -2249 125 -2227
rect 91 -2295 125 -2287
rect 91 -2321 125 -2295
rect 91 -2363 125 -2359
rect 91 -2393 125 -2363
rect 91 -2465 125 -2431
rect 199 2431 233 2465
rect 199 2363 233 2393
rect 199 2359 233 2363
rect 199 2295 233 2321
rect 199 2287 233 2295
rect 199 2227 233 2249
rect 199 2215 233 2227
rect 199 2159 233 2177
rect 199 2143 233 2159
rect 199 2091 233 2105
rect 199 2071 233 2091
rect 199 2023 233 2033
rect 199 1999 233 2023
rect 199 1955 233 1961
rect 199 1927 233 1955
rect 199 1887 233 1889
rect 199 1855 233 1887
rect 199 1785 233 1817
rect 199 1783 233 1785
rect 199 1717 233 1745
rect 199 1711 233 1717
rect 199 1649 233 1673
rect 199 1639 233 1649
rect 199 1581 233 1601
rect 199 1567 233 1581
rect 199 1513 233 1529
rect 199 1495 233 1513
rect 199 1445 233 1457
rect 199 1423 233 1445
rect 199 1377 233 1385
rect 199 1351 233 1377
rect 199 1309 233 1313
rect 199 1279 233 1309
rect 199 1207 233 1241
rect 199 1139 233 1169
rect 199 1135 233 1139
rect 199 1071 233 1097
rect 199 1063 233 1071
rect 199 1003 233 1025
rect 199 991 233 1003
rect 199 935 233 953
rect 199 919 233 935
rect 199 867 233 881
rect 199 847 233 867
rect 199 799 233 809
rect 199 775 233 799
rect 199 731 233 737
rect 199 703 233 731
rect 199 663 233 665
rect 199 631 233 663
rect 199 561 233 593
rect 199 559 233 561
rect 199 493 233 521
rect 199 487 233 493
rect 199 425 233 449
rect 199 415 233 425
rect 199 357 233 377
rect 199 343 233 357
rect 199 289 233 305
rect 199 271 233 289
rect 199 221 233 233
rect 199 199 233 221
rect 199 153 233 161
rect 199 127 233 153
rect 199 85 233 89
rect 199 55 233 85
rect 199 -17 233 17
rect 199 -85 233 -55
rect 199 -89 233 -85
rect 199 -153 233 -127
rect 199 -161 233 -153
rect 199 -221 233 -199
rect 199 -233 233 -221
rect 199 -289 233 -271
rect 199 -305 233 -289
rect 199 -357 233 -343
rect 199 -377 233 -357
rect 199 -425 233 -415
rect 199 -449 233 -425
rect 199 -493 233 -487
rect 199 -521 233 -493
rect 199 -561 233 -559
rect 199 -593 233 -561
rect 199 -663 233 -631
rect 199 -665 233 -663
rect 199 -731 233 -703
rect 199 -737 233 -731
rect 199 -799 233 -775
rect 199 -809 233 -799
rect 199 -867 233 -847
rect 199 -881 233 -867
rect 199 -935 233 -919
rect 199 -953 233 -935
rect 199 -1003 233 -991
rect 199 -1025 233 -1003
rect 199 -1071 233 -1063
rect 199 -1097 233 -1071
rect 199 -1139 233 -1135
rect 199 -1169 233 -1139
rect 199 -1241 233 -1207
rect 199 -1309 233 -1279
rect 199 -1313 233 -1309
rect 199 -1377 233 -1351
rect 199 -1385 233 -1377
rect 199 -1445 233 -1423
rect 199 -1457 233 -1445
rect 199 -1513 233 -1495
rect 199 -1529 233 -1513
rect 199 -1581 233 -1567
rect 199 -1601 233 -1581
rect 199 -1649 233 -1639
rect 199 -1673 233 -1649
rect 199 -1717 233 -1711
rect 199 -1745 233 -1717
rect 199 -1785 233 -1783
rect 199 -1817 233 -1785
rect 199 -1887 233 -1855
rect 199 -1889 233 -1887
rect 199 -1955 233 -1927
rect 199 -1961 233 -1955
rect 199 -2023 233 -1999
rect 199 -2033 233 -2023
rect 199 -2091 233 -2071
rect 199 -2105 233 -2091
rect 199 -2159 233 -2143
rect 199 -2177 233 -2159
rect 199 -2227 233 -2215
rect 199 -2249 233 -2227
rect 199 -2295 233 -2287
rect 199 -2321 233 -2295
rect 199 -2363 233 -2359
rect 199 -2393 233 -2363
rect 199 -2465 233 -2431
rect 307 2431 341 2465
rect 307 2363 341 2393
rect 307 2359 341 2363
rect 307 2295 341 2321
rect 307 2287 341 2295
rect 307 2227 341 2249
rect 307 2215 341 2227
rect 307 2159 341 2177
rect 307 2143 341 2159
rect 307 2091 341 2105
rect 307 2071 341 2091
rect 307 2023 341 2033
rect 307 1999 341 2023
rect 307 1955 341 1961
rect 307 1927 341 1955
rect 307 1887 341 1889
rect 307 1855 341 1887
rect 307 1785 341 1817
rect 307 1783 341 1785
rect 307 1717 341 1745
rect 307 1711 341 1717
rect 307 1649 341 1673
rect 307 1639 341 1649
rect 307 1581 341 1601
rect 307 1567 341 1581
rect 307 1513 341 1529
rect 307 1495 341 1513
rect 307 1445 341 1457
rect 307 1423 341 1445
rect 307 1377 341 1385
rect 307 1351 341 1377
rect 307 1309 341 1313
rect 307 1279 341 1309
rect 307 1207 341 1241
rect 307 1139 341 1169
rect 307 1135 341 1139
rect 307 1071 341 1097
rect 307 1063 341 1071
rect 307 1003 341 1025
rect 307 991 341 1003
rect 307 935 341 953
rect 307 919 341 935
rect 307 867 341 881
rect 307 847 341 867
rect 307 799 341 809
rect 307 775 341 799
rect 307 731 341 737
rect 307 703 341 731
rect 307 663 341 665
rect 307 631 341 663
rect 307 561 341 593
rect 307 559 341 561
rect 307 493 341 521
rect 307 487 341 493
rect 307 425 341 449
rect 307 415 341 425
rect 307 357 341 377
rect 307 343 341 357
rect 307 289 341 305
rect 307 271 341 289
rect 307 221 341 233
rect 307 199 341 221
rect 307 153 341 161
rect 307 127 341 153
rect 307 85 341 89
rect 307 55 341 85
rect 307 -17 341 17
rect 307 -85 341 -55
rect 307 -89 341 -85
rect 307 -153 341 -127
rect 307 -161 341 -153
rect 307 -221 341 -199
rect 307 -233 341 -221
rect 307 -289 341 -271
rect 307 -305 341 -289
rect 307 -357 341 -343
rect 307 -377 341 -357
rect 307 -425 341 -415
rect 307 -449 341 -425
rect 307 -493 341 -487
rect 307 -521 341 -493
rect 307 -561 341 -559
rect 307 -593 341 -561
rect 307 -663 341 -631
rect 307 -665 341 -663
rect 307 -731 341 -703
rect 307 -737 341 -731
rect 307 -799 341 -775
rect 307 -809 341 -799
rect 307 -867 341 -847
rect 307 -881 341 -867
rect 307 -935 341 -919
rect 307 -953 341 -935
rect 307 -1003 341 -991
rect 307 -1025 341 -1003
rect 307 -1071 341 -1063
rect 307 -1097 341 -1071
rect 307 -1139 341 -1135
rect 307 -1169 341 -1139
rect 307 -1241 341 -1207
rect 307 -1309 341 -1279
rect 307 -1313 341 -1309
rect 307 -1377 341 -1351
rect 307 -1385 341 -1377
rect 307 -1445 341 -1423
rect 307 -1457 341 -1445
rect 307 -1513 341 -1495
rect 307 -1529 341 -1513
rect 307 -1581 341 -1567
rect 307 -1601 341 -1581
rect 307 -1649 341 -1639
rect 307 -1673 341 -1649
rect 307 -1717 341 -1711
rect 307 -1745 341 -1717
rect 307 -1785 341 -1783
rect 307 -1817 341 -1785
rect 307 -1887 341 -1855
rect 307 -1889 341 -1887
rect 307 -1955 341 -1927
rect 307 -1961 341 -1955
rect 307 -2023 341 -1999
rect 307 -2033 341 -2023
rect 307 -2091 341 -2071
rect 307 -2105 341 -2091
rect 307 -2159 341 -2143
rect 307 -2177 341 -2159
rect 307 -2227 341 -2215
rect 307 -2249 341 -2227
rect 307 -2295 341 -2287
rect 307 -2321 341 -2295
rect 307 -2363 341 -2359
rect 307 -2393 341 -2363
rect 307 -2465 341 -2431
rect 415 2431 449 2465
rect 415 2363 449 2393
rect 415 2359 449 2363
rect 415 2295 449 2321
rect 415 2287 449 2295
rect 415 2227 449 2249
rect 415 2215 449 2227
rect 415 2159 449 2177
rect 415 2143 449 2159
rect 415 2091 449 2105
rect 415 2071 449 2091
rect 415 2023 449 2033
rect 415 1999 449 2023
rect 415 1955 449 1961
rect 415 1927 449 1955
rect 415 1887 449 1889
rect 415 1855 449 1887
rect 415 1785 449 1817
rect 415 1783 449 1785
rect 415 1717 449 1745
rect 415 1711 449 1717
rect 415 1649 449 1673
rect 415 1639 449 1649
rect 415 1581 449 1601
rect 415 1567 449 1581
rect 415 1513 449 1529
rect 415 1495 449 1513
rect 415 1445 449 1457
rect 415 1423 449 1445
rect 415 1377 449 1385
rect 415 1351 449 1377
rect 415 1309 449 1313
rect 415 1279 449 1309
rect 415 1207 449 1241
rect 415 1139 449 1169
rect 415 1135 449 1139
rect 415 1071 449 1097
rect 415 1063 449 1071
rect 415 1003 449 1025
rect 415 991 449 1003
rect 415 935 449 953
rect 415 919 449 935
rect 415 867 449 881
rect 415 847 449 867
rect 415 799 449 809
rect 415 775 449 799
rect 415 731 449 737
rect 415 703 449 731
rect 415 663 449 665
rect 415 631 449 663
rect 415 561 449 593
rect 415 559 449 561
rect 415 493 449 521
rect 415 487 449 493
rect 415 425 449 449
rect 415 415 449 425
rect 415 357 449 377
rect 415 343 449 357
rect 415 289 449 305
rect 415 271 449 289
rect 415 221 449 233
rect 415 199 449 221
rect 415 153 449 161
rect 415 127 449 153
rect 415 85 449 89
rect 415 55 449 85
rect 415 -17 449 17
rect 415 -85 449 -55
rect 415 -89 449 -85
rect 415 -153 449 -127
rect 415 -161 449 -153
rect 415 -221 449 -199
rect 415 -233 449 -221
rect 415 -289 449 -271
rect 415 -305 449 -289
rect 415 -357 449 -343
rect 415 -377 449 -357
rect 415 -425 449 -415
rect 415 -449 449 -425
rect 415 -493 449 -487
rect 415 -521 449 -493
rect 415 -561 449 -559
rect 415 -593 449 -561
rect 415 -663 449 -631
rect 415 -665 449 -663
rect 415 -731 449 -703
rect 415 -737 449 -731
rect 415 -799 449 -775
rect 415 -809 449 -799
rect 415 -867 449 -847
rect 415 -881 449 -867
rect 415 -935 449 -919
rect 415 -953 449 -935
rect 415 -1003 449 -991
rect 415 -1025 449 -1003
rect 415 -1071 449 -1063
rect 415 -1097 449 -1071
rect 415 -1139 449 -1135
rect 415 -1169 449 -1139
rect 415 -1241 449 -1207
rect 415 -1309 449 -1279
rect 415 -1313 449 -1309
rect 415 -1377 449 -1351
rect 415 -1385 449 -1377
rect 415 -1445 449 -1423
rect 415 -1457 449 -1445
rect 415 -1513 449 -1495
rect 415 -1529 449 -1513
rect 415 -1581 449 -1567
rect 415 -1601 449 -1581
rect 415 -1649 449 -1639
rect 415 -1673 449 -1649
rect 415 -1717 449 -1711
rect 415 -1745 449 -1717
rect 415 -1785 449 -1783
rect 415 -1817 449 -1785
rect 415 -1887 449 -1855
rect 415 -1889 449 -1887
rect 415 -1955 449 -1927
rect 415 -1961 449 -1955
rect 415 -2023 449 -1999
rect 415 -2033 449 -2023
rect 415 -2091 449 -2071
rect 415 -2105 449 -2091
rect 415 -2159 449 -2143
rect 415 -2177 449 -2159
rect 415 -2227 449 -2215
rect 415 -2249 449 -2227
rect 415 -2295 449 -2287
rect 415 -2321 449 -2295
rect 415 -2363 449 -2359
rect 415 -2393 449 -2363
rect 415 -2465 449 -2431
rect -395 -2581 -361 -2547
rect -179 -2581 -145 -2547
rect 37 -2581 71 -2547
rect 253 -2581 287 -2547
<< metal1 >>
rect -299 2581 -241 2587
rect -299 2547 -287 2581
rect -253 2547 -241 2581
rect -299 2541 -241 2547
rect -83 2581 -25 2587
rect -83 2547 -71 2581
rect -37 2547 -25 2581
rect -83 2541 -25 2547
rect 133 2581 191 2587
rect 133 2547 145 2581
rect 179 2547 191 2581
rect 133 2541 191 2547
rect 349 2581 407 2587
rect 349 2547 361 2581
rect 395 2547 407 2581
rect 349 2541 407 2547
rect -455 2465 -409 2500
rect -455 2431 -449 2465
rect -415 2431 -409 2465
rect -455 2393 -409 2431
rect -455 2359 -449 2393
rect -415 2359 -409 2393
rect -455 2321 -409 2359
rect -455 2287 -449 2321
rect -415 2287 -409 2321
rect -455 2249 -409 2287
rect -455 2215 -449 2249
rect -415 2215 -409 2249
rect -455 2177 -409 2215
rect -455 2143 -449 2177
rect -415 2143 -409 2177
rect -455 2105 -409 2143
rect -455 2071 -449 2105
rect -415 2071 -409 2105
rect -455 2033 -409 2071
rect -455 1999 -449 2033
rect -415 1999 -409 2033
rect -455 1961 -409 1999
rect -455 1927 -449 1961
rect -415 1927 -409 1961
rect -455 1889 -409 1927
rect -455 1855 -449 1889
rect -415 1855 -409 1889
rect -455 1817 -409 1855
rect -455 1783 -449 1817
rect -415 1783 -409 1817
rect -455 1745 -409 1783
rect -455 1711 -449 1745
rect -415 1711 -409 1745
rect -455 1673 -409 1711
rect -455 1639 -449 1673
rect -415 1639 -409 1673
rect -455 1601 -409 1639
rect -455 1567 -449 1601
rect -415 1567 -409 1601
rect -455 1529 -409 1567
rect -455 1495 -449 1529
rect -415 1495 -409 1529
rect -455 1457 -409 1495
rect -455 1423 -449 1457
rect -415 1423 -409 1457
rect -455 1385 -409 1423
rect -455 1351 -449 1385
rect -415 1351 -409 1385
rect -455 1313 -409 1351
rect -455 1279 -449 1313
rect -415 1279 -409 1313
rect -455 1241 -409 1279
rect -455 1207 -449 1241
rect -415 1207 -409 1241
rect -455 1169 -409 1207
rect -455 1135 -449 1169
rect -415 1135 -409 1169
rect -455 1097 -409 1135
rect -455 1063 -449 1097
rect -415 1063 -409 1097
rect -455 1025 -409 1063
rect -455 991 -449 1025
rect -415 991 -409 1025
rect -455 953 -409 991
rect -455 919 -449 953
rect -415 919 -409 953
rect -455 881 -409 919
rect -455 847 -449 881
rect -415 847 -409 881
rect -455 809 -409 847
rect -455 775 -449 809
rect -415 775 -409 809
rect -455 737 -409 775
rect -455 703 -449 737
rect -415 703 -409 737
rect -455 665 -409 703
rect -455 631 -449 665
rect -415 631 -409 665
rect -455 593 -409 631
rect -455 559 -449 593
rect -415 559 -409 593
rect -455 521 -409 559
rect -455 487 -449 521
rect -415 487 -409 521
rect -455 449 -409 487
rect -455 415 -449 449
rect -415 415 -409 449
rect -455 377 -409 415
rect -455 343 -449 377
rect -415 343 -409 377
rect -455 305 -409 343
rect -455 271 -449 305
rect -415 271 -409 305
rect -455 233 -409 271
rect -455 199 -449 233
rect -415 199 -409 233
rect -455 161 -409 199
rect -455 127 -449 161
rect -415 127 -409 161
rect -455 89 -409 127
rect -455 55 -449 89
rect -415 55 -409 89
rect -455 17 -409 55
rect -455 -17 -449 17
rect -415 -17 -409 17
rect -455 -55 -409 -17
rect -455 -89 -449 -55
rect -415 -89 -409 -55
rect -455 -127 -409 -89
rect -455 -161 -449 -127
rect -415 -161 -409 -127
rect -455 -199 -409 -161
rect -455 -233 -449 -199
rect -415 -233 -409 -199
rect -455 -271 -409 -233
rect -455 -305 -449 -271
rect -415 -305 -409 -271
rect -455 -343 -409 -305
rect -455 -377 -449 -343
rect -415 -377 -409 -343
rect -455 -415 -409 -377
rect -455 -449 -449 -415
rect -415 -449 -409 -415
rect -455 -487 -409 -449
rect -455 -521 -449 -487
rect -415 -521 -409 -487
rect -455 -559 -409 -521
rect -455 -593 -449 -559
rect -415 -593 -409 -559
rect -455 -631 -409 -593
rect -455 -665 -449 -631
rect -415 -665 -409 -631
rect -455 -703 -409 -665
rect -455 -737 -449 -703
rect -415 -737 -409 -703
rect -455 -775 -409 -737
rect -455 -809 -449 -775
rect -415 -809 -409 -775
rect -455 -847 -409 -809
rect -455 -881 -449 -847
rect -415 -881 -409 -847
rect -455 -919 -409 -881
rect -455 -953 -449 -919
rect -415 -953 -409 -919
rect -455 -991 -409 -953
rect -455 -1025 -449 -991
rect -415 -1025 -409 -991
rect -455 -1063 -409 -1025
rect -455 -1097 -449 -1063
rect -415 -1097 -409 -1063
rect -455 -1135 -409 -1097
rect -455 -1169 -449 -1135
rect -415 -1169 -409 -1135
rect -455 -1207 -409 -1169
rect -455 -1241 -449 -1207
rect -415 -1241 -409 -1207
rect -455 -1279 -409 -1241
rect -455 -1313 -449 -1279
rect -415 -1313 -409 -1279
rect -455 -1351 -409 -1313
rect -455 -1385 -449 -1351
rect -415 -1385 -409 -1351
rect -455 -1423 -409 -1385
rect -455 -1457 -449 -1423
rect -415 -1457 -409 -1423
rect -455 -1495 -409 -1457
rect -455 -1529 -449 -1495
rect -415 -1529 -409 -1495
rect -455 -1567 -409 -1529
rect -455 -1601 -449 -1567
rect -415 -1601 -409 -1567
rect -455 -1639 -409 -1601
rect -455 -1673 -449 -1639
rect -415 -1673 -409 -1639
rect -455 -1711 -409 -1673
rect -455 -1745 -449 -1711
rect -415 -1745 -409 -1711
rect -455 -1783 -409 -1745
rect -455 -1817 -449 -1783
rect -415 -1817 -409 -1783
rect -455 -1855 -409 -1817
rect -455 -1889 -449 -1855
rect -415 -1889 -409 -1855
rect -455 -1927 -409 -1889
rect -455 -1961 -449 -1927
rect -415 -1961 -409 -1927
rect -455 -1999 -409 -1961
rect -455 -2033 -449 -1999
rect -415 -2033 -409 -1999
rect -455 -2071 -409 -2033
rect -455 -2105 -449 -2071
rect -415 -2105 -409 -2071
rect -455 -2143 -409 -2105
rect -455 -2177 -449 -2143
rect -415 -2177 -409 -2143
rect -455 -2215 -409 -2177
rect -455 -2249 -449 -2215
rect -415 -2249 -409 -2215
rect -455 -2287 -409 -2249
rect -455 -2321 -449 -2287
rect -415 -2321 -409 -2287
rect -455 -2359 -409 -2321
rect -455 -2393 -449 -2359
rect -415 -2393 -409 -2359
rect -455 -2431 -409 -2393
rect -455 -2465 -449 -2431
rect -415 -2465 -409 -2431
rect -455 -2500 -409 -2465
rect -347 2465 -301 2500
rect -347 2431 -341 2465
rect -307 2431 -301 2465
rect -347 2393 -301 2431
rect -347 2359 -341 2393
rect -307 2359 -301 2393
rect -347 2321 -301 2359
rect -347 2287 -341 2321
rect -307 2287 -301 2321
rect -347 2249 -301 2287
rect -347 2215 -341 2249
rect -307 2215 -301 2249
rect -347 2177 -301 2215
rect -347 2143 -341 2177
rect -307 2143 -301 2177
rect -347 2105 -301 2143
rect -347 2071 -341 2105
rect -307 2071 -301 2105
rect -347 2033 -301 2071
rect -347 1999 -341 2033
rect -307 1999 -301 2033
rect -347 1961 -301 1999
rect -347 1927 -341 1961
rect -307 1927 -301 1961
rect -347 1889 -301 1927
rect -347 1855 -341 1889
rect -307 1855 -301 1889
rect -347 1817 -301 1855
rect -347 1783 -341 1817
rect -307 1783 -301 1817
rect -347 1745 -301 1783
rect -347 1711 -341 1745
rect -307 1711 -301 1745
rect -347 1673 -301 1711
rect -347 1639 -341 1673
rect -307 1639 -301 1673
rect -347 1601 -301 1639
rect -347 1567 -341 1601
rect -307 1567 -301 1601
rect -347 1529 -301 1567
rect -347 1495 -341 1529
rect -307 1495 -301 1529
rect -347 1457 -301 1495
rect -347 1423 -341 1457
rect -307 1423 -301 1457
rect -347 1385 -301 1423
rect -347 1351 -341 1385
rect -307 1351 -301 1385
rect -347 1313 -301 1351
rect -347 1279 -341 1313
rect -307 1279 -301 1313
rect -347 1241 -301 1279
rect -347 1207 -341 1241
rect -307 1207 -301 1241
rect -347 1169 -301 1207
rect -347 1135 -341 1169
rect -307 1135 -301 1169
rect -347 1097 -301 1135
rect -347 1063 -341 1097
rect -307 1063 -301 1097
rect -347 1025 -301 1063
rect -347 991 -341 1025
rect -307 991 -301 1025
rect -347 953 -301 991
rect -347 919 -341 953
rect -307 919 -301 953
rect -347 881 -301 919
rect -347 847 -341 881
rect -307 847 -301 881
rect -347 809 -301 847
rect -347 775 -341 809
rect -307 775 -301 809
rect -347 737 -301 775
rect -347 703 -341 737
rect -307 703 -301 737
rect -347 665 -301 703
rect -347 631 -341 665
rect -307 631 -301 665
rect -347 593 -301 631
rect -347 559 -341 593
rect -307 559 -301 593
rect -347 521 -301 559
rect -347 487 -341 521
rect -307 487 -301 521
rect -347 449 -301 487
rect -347 415 -341 449
rect -307 415 -301 449
rect -347 377 -301 415
rect -347 343 -341 377
rect -307 343 -301 377
rect -347 305 -301 343
rect -347 271 -341 305
rect -307 271 -301 305
rect -347 233 -301 271
rect -347 199 -341 233
rect -307 199 -301 233
rect -347 161 -301 199
rect -347 127 -341 161
rect -307 127 -301 161
rect -347 89 -301 127
rect -347 55 -341 89
rect -307 55 -301 89
rect -347 17 -301 55
rect -347 -17 -341 17
rect -307 -17 -301 17
rect -347 -55 -301 -17
rect -347 -89 -341 -55
rect -307 -89 -301 -55
rect -347 -127 -301 -89
rect -347 -161 -341 -127
rect -307 -161 -301 -127
rect -347 -199 -301 -161
rect -347 -233 -341 -199
rect -307 -233 -301 -199
rect -347 -271 -301 -233
rect -347 -305 -341 -271
rect -307 -305 -301 -271
rect -347 -343 -301 -305
rect -347 -377 -341 -343
rect -307 -377 -301 -343
rect -347 -415 -301 -377
rect -347 -449 -341 -415
rect -307 -449 -301 -415
rect -347 -487 -301 -449
rect -347 -521 -341 -487
rect -307 -521 -301 -487
rect -347 -559 -301 -521
rect -347 -593 -341 -559
rect -307 -593 -301 -559
rect -347 -631 -301 -593
rect -347 -665 -341 -631
rect -307 -665 -301 -631
rect -347 -703 -301 -665
rect -347 -737 -341 -703
rect -307 -737 -301 -703
rect -347 -775 -301 -737
rect -347 -809 -341 -775
rect -307 -809 -301 -775
rect -347 -847 -301 -809
rect -347 -881 -341 -847
rect -307 -881 -301 -847
rect -347 -919 -301 -881
rect -347 -953 -341 -919
rect -307 -953 -301 -919
rect -347 -991 -301 -953
rect -347 -1025 -341 -991
rect -307 -1025 -301 -991
rect -347 -1063 -301 -1025
rect -347 -1097 -341 -1063
rect -307 -1097 -301 -1063
rect -347 -1135 -301 -1097
rect -347 -1169 -341 -1135
rect -307 -1169 -301 -1135
rect -347 -1207 -301 -1169
rect -347 -1241 -341 -1207
rect -307 -1241 -301 -1207
rect -347 -1279 -301 -1241
rect -347 -1313 -341 -1279
rect -307 -1313 -301 -1279
rect -347 -1351 -301 -1313
rect -347 -1385 -341 -1351
rect -307 -1385 -301 -1351
rect -347 -1423 -301 -1385
rect -347 -1457 -341 -1423
rect -307 -1457 -301 -1423
rect -347 -1495 -301 -1457
rect -347 -1529 -341 -1495
rect -307 -1529 -301 -1495
rect -347 -1567 -301 -1529
rect -347 -1601 -341 -1567
rect -307 -1601 -301 -1567
rect -347 -1639 -301 -1601
rect -347 -1673 -341 -1639
rect -307 -1673 -301 -1639
rect -347 -1711 -301 -1673
rect -347 -1745 -341 -1711
rect -307 -1745 -301 -1711
rect -347 -1783 -301 -1745
rect -347 -1817 -341 -1783
rect -307 -1817 -301 -1783
rect -347 -1855 -301 -1817
rect -347 -1889 -341 -1855
rect -307 -1889 -301 -1855
rect -347 -1927 -301 -1889
rect -347 -1961 -341 -1927
rect -307 -1961 -301 -1927
rect -347 -1999 -301 -1961
rect -347 -2033 -341 -1999
rect -307 -2033 -301 -1999
rect -347 -2071 -301 -2033
rect -347 -2105 -341 -2071
rect -307 -2105 -301 -2071
rect -347 -2143 -301 -2105
rect -347 -2177 -341 -2143
rect -307 -2177 -301 -2143
rect -347 -2215 -301 -2177
rect -347 -2249 -341 -2215
rect -307 -2249 -301 -2215
rect -347 -2287 -301 -2249
rect -347 -2321 -341 -2287
rect -307 -2321 -301 -2287
rect -347 -2359 -301 -2321
rect -347 -2393 -341 -2359
rect -307 -2393 -301 -2359
rect -347 -2431 -301 -2393
rect -347 -2465 -341 -2431
rect -307 -2465 -301 -2431
rect -347 -2500 -301 -2465
rect -239 2465 -193 2500
rect -239 2431 -233 2465
rect -199 2431 -193 2465
rect -239 2393 -193 2431
rect -239 2359 -233 2393
rect -199 2359 -193 2393
rect -239 2321 -193 2359
rect -239 2287 -233 2321
rect -199 2287 -193 2321
rect -239 2249 -193 2287
rect -239 2215 -233 2249
rect -199 2215 -193 2249
rect -239 2177 -193 2215
rect -239 2143 -233 2177
rect -199 2143 -193 2177
rect -239 2105 -193 2143
rect -239 2071 -233 2105
rect -199 2071 -193 2105
rect -239 2033 -193 2071
rect -239 1999 -233 2033
rect -199 1999 -193 2033
rect -239 1961 -193 1999
rect -239 1927 -233 1961
rect -199 1927 -193 1961
rect -239 1889 -193 1927
rect -239 1855 -233 1889
rect -199 1855 -193 1889
rect -239 1817 -193 1855
rect -239 1783 -233 1817
rect -199 1783 -193 1817
rect -239 1745 -193 1783
rect -239 1711 -233 1745
rect -199 1711 -193 1745
rect -239 1673 -193 1711
rect -239 1639 -233 1673
rect -199 1639 -193 1673
rect -239 1601 -193 1639
rect -239 1567 -233 1601
rect -199 1567 -193 1601
rect -239 1529 -193 1567
rect -239 1495 -233 1529
rect -199 1495 -193 1529
rect -239 1457 -193 1495
rect -239 1423 -233 1457
rect -199 1423 -193 1457
rect -239 1385 -193 1423
rect -239 1351 -233 1385
rect -199 1351 -193 1385
rect -239 1313 -193 1351
rect -239 1279 -233 1313
rect -199 1279 -193 1313
rect -239 1241 -193 1279
rect -239 1207 -233 1241
rect -199 1207 -193 1241
rect -239 1169 -193 1207
rect -239 1135 -233 1169
rect -199 1135 -193 1169
rect -239 1097 -193 1135
rect -239 1063 -233 1097
rect -199 1063 -193 1097
rect -239 1025 -193 1063
rect -239 991 -233 1025
rect -199 991 -193 1025
rect -239 953 -193 991
rect -239 919 -233 953
rect -199 919 -193 953
rect -239 881 -193 919
rect -239 847 -233 881
rect -199 847 -193 881
rect -239 809 -193 847
rect -239 775 -233 809
rect -199 775 -193 809
rect -239 737 -193 775
rect -239 703 -233 737
rect -199 703 -193 737
rect -239 665 -193 703
rect -239 631 -233 665
rect -199 631 -193 665
rect -239 593 -193 631
rect -239 559 -233 593
rect -199 559 -193 593
rect -239 521 -193 559
rect -239 487 -233 521
rect -199 487 -193 521
rect -239 449 -193 487
rect -239 415 -233 449
rect -199 415 -193 449
rect -239 377 -193 415
rect -239 343 -233 377
rect -199 343 -193 377
rect -239 305 -193 343
rect -239 271 -233 305
rect -199 271 -193 305
rect -239 233 -193 271
rect -239 199 -233 233
rect -199 199 -193 233
rect -239 161 -193 199
rect -239 127 -233 161
rect -199 127 -193 161
rect -239 89 -193 127
rect -239 55 -233 89
rect -199 55 -193 89
rect -239 17 -193 55
rect -239 -17 -233 17
rect -199 -17 -193 17
rect -239 -55 -193 -17
rect -239 -89 -233 -55
rect -199 -89 -193 -55
rect -239 -127 -193 -89
rect -239 -161 -233 -127
rect -199 -161 -193 -127
rect -239 -199 -193 -161
rect -239 -233 -233 -199
rect -199 -233 -193 -199
rect -239 -271 -193 -233
rect -239 -305 -233 -271
rect -199 -305 -193 -271
rect -239 -343 -193 -305
rect -239 -377 -233 -343
rect -199 -377 -193 -343
rect -239 -415 -193 -377
rect -239 -449 -233 -415
rect -199 -449 -193 -415
rect -239 -487 -193 -449
rect -239 -521 -233 -487
rect -199 -521 -193 -487
rect -239 -559 -193 -521
rect -239 -593 -233 -559
rect -199 -593 -193 -559
rect -239 -631 -193 -593
rect -239 -665 -233 -631
rect -199 -665 -193 -631
rect -239 -703 -193 -665
rect -239 -737 -233 -703
rect -199 -737 -193 -703
rect -239 -775 -193 -737
rect -239 -809 -233 -775
rect -199 -809 -193 -775
rect -239 -847 -193 -809
rect -239 -881 -233 -847
rect -199 -881 -193 -847
rect -239 -919 -193 -881
rect -239 -953 -233 -919
rect -199 -953 -193 -919
rect -239 -991 -193 -953
rect -239 -1025 -233 -991
rect -199 -1025 -193 -991
rect -239 -1063 -193 -1025
rect -239 -1097 -233 -1063
rect -199 -1097 -193 -1063
rect -239 -1135 -193 -1097
rect -239 -1169 -233 -1135
rect -199 -1169 -193 -1135
rect -239 -1207 -193 -1169
rect -239 -1241 -233 -1207
rect -199 -1241 -193 -1207
rect -239 -1279 -193 -1241
rect -239 -1313 -233 -1279
rect -199 -1313 -193 -1279
rect -239 -1351 -193 -1313
rect -239 -1385 -233 -1351
rect -199 -1385 -193 -1351
rect -239 -1423 -193 -1385
rect -239 -1457 -233 -1423
rect -199 -1457 -193 -1423
rect -239 -1495 -193 -1457
rect -239 -1529 -233 -1495
rect -199 -1529 -193 -1495
rect -239 -1567 -193 -1529
rect -239 -1601 -233 -1567
rect -199 -1601 -193 -1567
rect -239 -1639 -193 -1601
rect -239 -1673 -233 -1639
rect -199 -1673 -193 -1639
rect -239 -1711 -193 -1673
rect -239 -1745 -233 -1711
rect -199 -1745 -193 -1711
rect -239 -1783 -193 -1745
rect -239 -1817 -233 -1783
rect -199 -1817 -193 -1783
rect -239 -1855 -193 -1817
rect -239 -1889 -233 -1855
rect -199 -1889 -193 -1855
rect -239 -1927 -193 -1889
rect -239 -1961 -233 -1927
rect -199 -1961 -193 -1927
rect -239 -1999 -193 -1961
rect -239 -2033 -233 -1999
rect -199 -2033 -193 -1999
rect -239 -2071 -193 -2033
rect -239 -2105 -233 -2071
rect -199 -2105 -193 -2071
rect -239 -2143 -193 -2105
rect -239 -2177 -233 -2143
rect -199 -2177 -193 -2143
rect -239 -2215 -193 -2177
rect -239 -2249 -233 -2215
rect -199 -2249 -193 -2215
rect -239 -2287 -193 -2249
rect -239 -2321 -233 -2287
rect -199 -2321 -193 -2287
rect -239 -2359 -193 -2321
rect -239 -2393 -233 -2359
rect -199 -2393 -193 -2359
rect -239 -2431 -193 -2393
rect -239 -2465 -233 -2431
rect -199 -2465 -193 -2431
rect -239 -2500 -193 -2465
rect -131 2465 -85 2500
rect -131 2431 -125 2465
rect -91 2431 -85 2465
rect -131 2393 -85 2431
rect -131 2359 -125 2393
rect -91 2359 -85 2393
rect -131 2321 -85 2359
rect -131 2287 -125 2321
rect -91 2287 -85 2321
rect -131 2249 -85 2287
rect -131 2215 -125 2249
rect -91 2215 -85 2249
rect -131 2177 -85 2215
rect -131 2143 -125 2177
rect -91 2143 -85 2177
rect -131 2105 -85 2143
rect -131 2071 -125 2105
rect -91 2071 -85 2105
rect -131 2033 -85 2071
rect -131 1999 -125 2033
rect -91 1999 -85 2033
rect -131 1961 -85 1999
rect -131 1927 -125 1961
rect -91 1927 -85 1961
rect -131 1889 -85 1927
rect -131 1855 -125 1889
rect -91 1855 -85 1889
rect -131 1817 -85 1855
rect -131 1783 -125 1817
rect -91 1783 -85 1817
rect -131 1745 -85 1783
rect -131 1711 -125 1745
rect -91 1711 -85 1745
rect -131 1673 -85 1711
rect -131 1639 -125 1673
rect -91 1639 -85 1673
rect -131 1601 -85 1639
rect -131 1567 -125 1601
rect -91 1567 -85 1601
rect -131 1529 -85 1567
rect -131 1495 -125 1529
rect -91 1495 -85 1529
rect -131 1457 -85 1495
rect -131 1423 -125 1457
rect -91 1423 -85 1457
rect -131 1385 -85 1423
rect -131 1351 -125 1385
rect -91 1351 -85 1385
rect -131 1313 -85 1351
rect -131 1279 -125 1313
rect -91 1279 -85 1313
rect -131 1241 -85 1279
rect -131 1207 -125 1241
rect -91 1207 -85 1241
rect -131 1169 -85 1207
rect -131 1135 -125 1169
rect -91 1135 -85 1169
rect -131 1097 -85 1135
rect -131 1063 -125 1097
rect -91 1063 -85 1097
rect -131 1025 -85 1063
rect -131 991 -125 1025
rect -91 991 -85 1025
rect -131 953 -85 991
rect -131 919 -125 953
rect -91 919 -85 953
rect -131 881 -85 919
rect -131 847 -125 881
rect -91 847 -85 881
rect -131 809 -85 847
rect -131 775 -125 809
rect -91 775 -85 809
rect -131 737 -85 775
rect -131 703 -125 737
rect -91 703 -85 737
rect -131 665 -85 703
rect -131 631 -125 665
rect -91 631 -85 665
rect -131 593 -85 631
rect -131 559 -125 593
rect -91 559 -85 593
rect -131 521 -85 559
rect -131 487 -125 521
rect -91 487 -85 521
rect -131 449 -85 487
rect -131 415 -125 449
rect -91 415 -85 449
rect -131 377 -85 415
rect -131 343 -125 377
rect -91 343 -85 377
rect -131 305 -85 343
rect -131 271 -125 305
rect -91 271 -85 305
rect -131 233 -85 271
rect -131 199 -125 233
rect -91 199 -85 233
rect -131 161 -85 199
rect -131 127 -125 161
rect -91 127 -85 161
rect -131 89 -85 127
rect -131 55 -125 89
rect -91 55 -85 89
rect -131 17 -85 55
rect -131 -17 -125 17
rect -91 -17 -85 17
rect -131 -55 -85 -17
rect -131 -89 -125 -55
rect -91 -89 -85 -55
rect -131 -127 -85 -89
rect -131 -161 -125 -127
rect -91 -161 -85 -127
rect -131 -199 -85 -161
rect -131 -233 -125 -199
rect -91 -233 -85 -199
rect -131 -271 -85 -233
rect -131 -305 -125 -271
rect -91 -305 -85 -271
rect -131 -343 -85 -305
rect -131 -377 -125 -343
rect -91 -377 -85 -343
rect -131 -415 -85 -377
rect -131 -449 -125 -415
rect -91 -449 -85 -415
rect -131 -487 -85 -449
rect -131 -521 -125 -487
rect -91 -521 -85 -487
rect -131 -559 -85 -521
rect -131 -593 -125 -559
rect -91 -593 -85 -559
rect -131 -631 -85 -593
rect -131 -665 -125 -631
rect -91 -665 -85 -631
rect -131 -703 -85 -665
rect -131 -737 -125 -703
rect -91 -737 -85 -703
rect -131 -775 -85 -737
rect -131 -809 -125 -775
rect -91 -809 -85 -775
rect -131 -847 -85 -809
rect -131 -881 -125 -847
rect -91 -881 -85 -847
rect -131 -919 -85 -881
rect -131 -953 -125 -919
rect -91 -953 -85 -919
rect -131 -991 -85 -953
rect -131 -1025 -125 -991
rect -91 -1025 -85 -991
rect -131 -1063 -85 -1025
rect -131 -1097 -125 -1063
rect -91 -1097 -85 -1063
rect -131 -1135 -85 -1097
rect -131 -1169 -125 -1135
rect -91 -1169 -85 -1135
rect -131 -1207 -85 -1169
rect -131 -1241 -125 -1207
rect -91 -1241 -85 -1207
rect -131 -1279 -85 -1241
rect -131 -1313 -125 -1279
rect -91 -1313 -85 -1279
rect -131 -1351 -85 -1313
rect -131 -1385 -125 -1351
rect -91 -1385 -85 -1351
rect -131 -1423 -85 -1385
rect -131 -1457 -125 -1423
rect -91 -1457 -85 -1423
rect -131 -1495 -85 -1457
rect -131 -1529 -125 -1495
rect -91 -1529 -85 -1495
rect -131 -1567 -85 -1529
rect -131 -1601 -125 -1567
rect -91 -1601 -85 -1567
rect -131 -1639 -85 -1601
rect -131 -1673 -125 -1639
rect -91 -1673 -85 -1639
rect -131 -1711 -85 -1673
rect -131 -1745 -125 -1711
rect -91 -1745 -85 -1711
rect -131 -1783 -85 -1745
rect -131 -1817 -125 -1783
rect -91 -1817 -85 -1783
rect -131 -1855 -85 -1817
rect -131 -1889 -125 -1855
rect -91 -1889 -85 -1855
rect -131 -1927 -85 -1889
rect -131 -1961 -125 -1927
rect -91 -1961 -85 -1927
rect -131 -1999 -85 -1961
rect -131 -2033 -125 -1999
rect -91 -2033 -85 -1999
rect -131 -2071 -85 -2033
rect -131 -2105 -125 -2071
rect -91 -2105 -85 -2071
rect -131 -2143 -85 -2105
rect -131 -2177 -125 -2143
rect -91 -2177 -85 -2143
rect -131 -2215 -85 -2177
rect -131 -2249 -125 -2215
rect -91 -2249 -85 -2215
rect -131 -2287 -85 -2249
rect -131 -2321 -125 -2287
rect -91 -2321 -85 -2287
rect -131 -2359 -85 -2321
rect -131 -2393 -125 -2359
rect -91 -2393 -85 -2359
rect -131 -2431 -85 -2393
rect -131 -2465 -125 -2431
rect -91 -2465 -85 -2431
rect -131 -2500 -85 -2465
rect -23 2465 23 2500
rect -23 2431 -17 2465
rect 17 2431 23 2465
rect -23 2393 23 2431
rect -23 2359 -17 2393
rect 17 2359 23 2393
rect -23 2321 23 2359
rect -23 2287 -17 2321
rect 17 2287 23 2321
rect -23 2249 23 2287
rect -23 2215 -17 2249
rect 17 2215 23 2249
rect -23 2177 23 2215
rect -23 2143 -17 2177
rect 17 2143 23 2177
rect -23 2105 23 2143
rect -23 2071 -17 2105
rect 17 2071 23 2105
rect -23 2033 23 2071
rect -23 1999 -17 2033
rect 17 1999 23 2033
rect -23 1961 23 1999
rect -23 1927 -17 1961
rect 17 1927 23 1961
rect -23 1889 23 1927
rect -23 1855 -17 1889
rect 17 1855 23 1889
rect -23 1817 23 1855
rect -23 1783 -17 1817
rect 17 1783 23 1817
rect -23 1745 23 1783
rect -23 1711 -17 1745
rect 17 1711 23 1745
rect -23 1673 23 1711
rect -23 1639 -17 1673
rect 17 1639 23 1673
rect -23 1601 23 1639
rect -23 1567 -17 1601
rect 17 1567 23 1601
rect -23 1529 23 1567
rect -23 1495 -17 1529
rect 17 1495 23 1529
rect -23 1457 23 1495
rect -23 1423 -17 1457
rect 17 1423 23 1457
rect -23 1385 23 1423
rect -23 1351 -17 1385
rect 17 1351 23 1385
rect -23 1313 23 1351
rect -23 1279 -17 1313
rect 17 1279 23 1313
rect -23 1241 23 1279
rect -23 1207 -17 1241
rect 17 1207 23 1241
rect -23 1169 23 1207
rect -23 1135 -17 1169
rect 17 1135 23 1169
rect -23 1097 23 1135
rect -23 1063 -17 1097
rect 17 1063 23 1097
rect -23 1025 23 1063
rect -23 991 -17 1025
rect 17 991 23 1025
rect -23 953 23 991
rect -23 919 -17 953
rect 17 919 23 953
rect -23 881 23 919
rect -23 847 -17 881
rect 17 847 23 881
rect -23 809 23 847
rect -23 775 -17 809
rect 17 775 23 809
rect -23 737 23 775
rect -23 703 -17 737
rect 17 703 23 737
rect -23 665 23 703
rect -23 631 -17 665
rect 17 631 23 665
rect -23 593 23 631
rect -23 559 -17 593
rect 17 559 23 593
rect -23 521 23 559
rect -23 487 -17 521
rect 17 487 23 521
rect -23 449 23 487
rect -23 415 -17 449
rect 17 415 23 449
rect -23 377 23 415
rect -23 343 -17 377
rect 17 343 23 377
rect -23 305 23 343
rect -23 271 -17 305
rect 17 271 23 305
rect -23 233 23 271
rect -23 199 -17 233
rect 17 199 23 233
rect -23 161 23 199
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -199 23 -161
rect -23 -233 -17 -199
rect 17 -233 23 -199
rect -23 -271 23 -233
rect -23 -305 -17 -271
rect 17 -305 23 -271
rect -23 -343 23 -305
rect -23 -377 -17 -343
rect 17 -377 23 -343
rect -23 -415 23 -377
rect -23 -449 -17 -415
rect 17 -449 23 -415
rect -23 -487 23 -449
rect -23 -521 -17 -487
rect 17 -521 23 -487
rect -23 -559 23 -521
rect -23 -593 -17 -559
rect 17 -593 23 -559
rect -23 -631 23 -593
rect -23 -665 -17 -631
rect 17 -665 23 -631
rect -23 -703 23 -665
rect -23 -737 -17 -703
rect 17 -737 23 -703
rect -23 -775 23 -737
rect -23 -809 -17 -775
rect 17 -809 23 -775
rect -23 -847 23 -809
rect -23 -881 -17 -847
rect 17 -881 23 -847
rect -23 -919 23 -881
rect -23 -953 -17 -919
rect 17 -953 23 -919
rect -23 -991 23 -953
rect -23 -1025 -17 -991
rect 17 -1025 23 -991
rect -23 -1063 23 -1025
rect -23 -1097 -17 -1063
rect 17 -1097 23 -1063
rect -23 -1135 23 -1097
rect -23 -1169 -17 -1135
rect 17 -1169 23 -1135
rect -23 -1207 23 -1169
rect -23 -1241 -17 -1207
rect 17 -1241 23 -1207
rect -23 -1279 23 -1241
rect -23 -1313 -17 -1279
rect 17 -1313 23 -1279
rect -23 -1351 23 -1313
rect -23 -1385 -17 -1351
rect 17 -1385 23 -1351
rect -23 -1423 23 -1385
rect -23 -1457 -17 -1423
rect 17 -1457 23 -1423
rect -23 -1495 23 -1457
rect -23 -1529 -17 -1495
rect 17 -1529 23 -1495
rect -23 -1567 23 -1529
rect -23 -1601 -17 -1567
rect 17 -1601 23 -1567
rect -23 -1639 23 -1601
rect -23 -1673 -17 -1639
rect 17 -1673 23 -1639
rect -23 -1711 23 -1673
rect -23 -1745 -17 -1711
rect 17 -1745 23 -1711
rect -23 -1783 23 -1745
rect -23 -1817 -17 -1783
rect 17 -1817 23 -1783
rect -23 -1855 23 -1817
rect -23 -1889 -17 -1855
rect 17 -1889 23 -1855
rect -23 -1927 23 -1889
rect -23 -1961 -17 -1927
rect 17 -1961 23 -1927
rect -23 -1999 23 -1961
rect -23 -2033 -17 -1999
rect 17 -2033 23 -1999
rect -23 -2071 23 -2033
rect -23 -2105 -17 -2071
rect 17 -2105 23 -2071
rect -23 -2143 23 -2105
rect -23 -2177 -17 -2143
rect 17 -2177 23 -2143
rect -23 -2215 23 -2177
rect -23 -2249 -17 -2215
rect 17 -2249 23 -2215
rect -23 -2287 23 -2249
rect -23 -2321 -17 -2287
rect 17 -2321 23 -2287
rect -23 -2359 23 -2321
rect -23 -2393 -17 -2359
rect 17 -2393 23 -2359
rect -23 -2431 23 -2393
rect -23 -2465 -17 -2431
rect 17 -2465 23 -2431
rect -23 -2500 23 -2465
rect 85 2465 131 2500
rect 85 2431 91 2465
rect 125 2431 131 2465
rect 85 2393 131 2431
rect 85 2359 91 2393
rect 125 2359 131 2393
rect 85 2321 131 2359
rect 85 2287 91 2321
rect 125 2287 131 2321
rect 85 2249 131 2287
rect 85 2215 91 2249
rect 125 2215 131 2249
rect 85 2177 131 2215
rect 85 2143 91 2177
rect 125 2143 131 2177
rect 85 2105 131 2143
rect 85 2071 91 2105
rect 125 2071 131 2105
rect 85 2033 131 2071
rect 85 1999 91 2033
rect 125 1999 131 2033
rect 85 1961 131 1999
rect 85 1927 91 1961
rect 125 1927 131 1961
rect 85 1889 131 1927
rect 85 1855 91 1889
rect 125 1855 131 1889
rect 85 1817 131 1855
rect 85 1783 91 1817
rect 125 1783 131 1817
rect 85 1745 131 1783
rect 85 1711 91 1745
rect 125 1711 131 1745
rect 85 1673 131 1711
rect 85 1639 91 1673
rect 125 1639 131 1673
rect 85 1601 131 1639
rect 85 1567 91 1601
rect 125 1567 131 1601
rect 85 1529 131 1567
rect 85 1495 91 1529
rect 125 1495 131 1529
rect 85 1457 131 1495
rect 85 1423 91 1457
rect 125 1423 131 1457
rect 85 1385 131 1423
rect 85 1351 91 1385
rect 125 1351 131 1385
rect 85 1313 131 1351
rect 85 1279 91 1313
rect 125 1279 131 1313
rect 85 1241 131 1279
rect 85 1207 91 1241
rect 125 1207 131 1241
rect 85 1169 131 1207
rect 85 1135 91 1169
rect 125 1135 131 1169
rect 85 1097 131 1135
rect 85 1063 91 1097
rect 125 1063 131 1097
rect 85 1025 131 1063
rect 85 991 91 1025
rect 125 991 131 1025
rect 85 953 131 991
rect 85 919 91 953
rect 125 919 131 953
rect 85 881 131 919
rect 85 847 91 881
rect 125 847 131 881
rect 85 809 131 847
rect 85 775 91 809
rect 125 775 131 809
rect 85 737 131 775
rect 85 703 91 737
rect 125 703 131 737
rect 85 665 131 703
rect 85 631 91 665
rect 125 631 131 665
rect 85 593 131 631
rect 85 559 91 593
rect 125 559 131 593
rect 85 521 131 559
rect 85 487 91 521
rect 125 487 131 521
rect 85 449 131 487
rect 85 415 91 449
rect 125 415 131 449
rect 85 377 131 415
rect 85 343 91 377
rect 125 343 131 377
rect 85 305 131 343
rect 85 271 91 305
rect 125 271 131 305
rect 85 233 131 271
rect 85 199 91 233
rect 125 199 131 233
rect 85 161 131 199
rect 85 127 91 161
rect 125 127 131 161
rect 85 89 131 127
rect 85 55 91 89
rect 125 55 131 89
rect 85 17 131 55
rect 85 -17 91 17
rect 125 -17 131 17
rect 85 -55 131 -17
rect 85 -89 91 -55
rect 125 -89 131 -55
rect 85 -127 131 -89
rect 85 -161 91 -127
rect 125 -161 131 -127
rect 85 -199 131 -161
rect 85 -233 91 -199
rect 125 -233 131 -199
rect 85 -271 131 -233
rect 85 -305 91 -271
rect 125 -305 131 -271
rect 85 -343 131 -305
rect 85 -377 91 -343
rect 125 -377 131 -343
rect 85 -415 131 -377
rect 85 -449 91 -415
rect 125 -449 131 -415
rect 85 -487 131 -449
rect 85 -521 91 -487
rect 125 -521 131 -487
rect 85 -559 131 -521
rect 85 -593 91 -559
rect 125 -593 131 -559
rect 85 -631 131 -593
rect 85 -665 91 -631
rect 125 -665 131 -631
rect 85 -703 131 -665
rect 85 -737 91 -703
rect 125 -737 131 -703
rect 85 -775 131 -737
rect 85 -809 91 -775
rect 125 -809 131 -775
rect 85 -847 131 -809
rect 85 -881 91 -847
rect 125 -881 131 -847
rect 85 -919 131 -881
rect 85 -953 91 -919
rect 125 -953 131 -919
rect 85 -991 131 -953
rect 85 -1025 91 -991
rect 125 -1025 131 -991
rect 85 -1063 131 -1025
rect 85 -1097 91 -1063
rect 125 -1097 131 -1063
rect 85 -1135 131 -1097
rect 85 -1169 91 -1135
rect 125 -1169 131 -1135
rect 85 -1207 131 -1169
rect 85 -1241 91 -1207
rect 125 -1241 131 -1207
rect 85 -1279 131 -1241
rect 85 -1313 91 -1279
rect 125 -1313 131 -1279
rect 85 -1351 131 -1313
rect 85 -1385 91 -1351
rect 125 -1385 131 -1351
rect 85 -1423 131 -1385
rect 85 -1457 91 -1423
rect 125 -1457 131 -1423
rect 85 -1495 131 -1457
rect 85 -1529 91 -1495
rect 125 -1529 131 -1495
rect 85 -1567 131 -1529
rect 85 -1601 91 -1567
rect 125 -1601 131 -1567
rect 85 -1639 131 -1601
rect 85 -1673 91 -1639
rect 125 -1673 131 -1639
rect 85 -1711 131 -1673
rect 85 -1745 91 -1711
rect 125 -1745 131 -1711
rect 85 -1783 131 -1745
rect 85 -1817 91 -1783
rect 125 -1817 131 -1783
rect 85 -1855 131 -1817
rect 85 -1889 91 -1855
rect 125 -1889 131 -1855
rect 85 -1927 131 -1889
rect 85 -1961 91 -1927
rect 125 -1961 131 -1927
rect 85 -1999 131 -1961
rect 85 -2033 91 -1999
rect 125 -2033 131 -1999
rect 85 -2071 131 -2033
rect 85 -2105 91 -2071
rect 125 -2105 131 -2071
rect 85 -2143 131 -2105
rect 85 -2177 91 -2143
rect 125 -2177 131 -2143
rect 85 -2215 131 -2177
rect 85 -2249 91 -2215
rect 125 -2249 131 -2215
rect 85 -2287 131 -2249
rect 85 -2321 91 -2287
rect 125 -2321 131 -2287
rect 85 -2359 131 -2321
rect 85 -2393 91 -2359
rect 125 -2393 131 -2359
rect 85 -2431 131 -2393
rect 85 -2465 91 -2431
rect 125 -2465 131 -2431
rect 85 -2500 131 -2465
rect 193 2465 239 2500
rect 193 2431 199 2465
rect 233 2431 239 2465
rect 193 2393 239 2431
rect 193 2359 199 2393
rect 233 2359 239 2393
rect 193 2321 239 2359
rect 193 2287 199 2321
rect 233 2287 239 2321
rect 193 2249 239 2287
rect 193 2215 199 2249
rect 233 2215 239 2249
rect 193 2177 239 2215
rect 193 2143 199 2177
rect 233 2143 239 2177
rect 193 2105 239 2143
rect 193 2071 199 2105
rect 233 2071 239 2105
rect 193 2033 239 2071
rect 193 1999 199 2033
rect 233 1999 239 2033
rect 193 1961 239 1999
rect 193 1927 199 1961
rect 233 1927 239 1961
rect 193 1889 239 1927
rect 193 1855 199 1889
rect 233 1855 239 1889
rect 193 1817 239 1855
rect 193 1783 199 1817
rect 233 1783 239 1817
rect 193 1745 239 1783
rect 193 1711 199 1745
rect 233 1711 239 1745
rect 193 1673 239 1711
rect 193 1639 199 1673
rect 233 1639 239 1673
rect 193 1601 239 1639
rect 193 1567 199 1601
rect 233 1567 239 1601
rect 193 1529 239 1567
rect 193 1495 199 1529
rect 233 1495 239 1529
rect 193 1457 239 1495
rect 193 1423 199 1457
rect 233 1423 239 1457
rect 193 1385 239 1423
rect 193 1351 199 1385
rect 233 1351 239 1385
rect 193 1313 239 1351
rect 193 1279 199 1313
rect 233 1279 239 1313
rect 193 1241 239 1279
rect 193 1207 199 1241
rect 233 1207 239 1241
rect 193 1169 239 1207
rect 193 1135 199 1169
rect 233 1135 239 1169
rect 193 1097 239 1135
rect 193 1063 199 1097
rect 233 1063 239 1097
rect 193 1025 239 1063
rect 193 991 199 1025
rect 233 991 239 1025
rect 193 953 239 991
rect 193 919 199 953
rect 233 919 239 953
rect 193 881 239 919
rect 193 847 199 881
rect 233 847 239 881
rect 193 809 239 847
rect 193 775 199 809
rect 233 775 239 809
rect 193 737 239 775
rect 193 703 199 737
rect 233 703 239 737
rect 193 665 239 703
rect 193 631 199 665
rect 233 631 239 665
rect 193 593 239 631
rect 193 559 199 593
rect 233 559 239 593
rect 193 521 239 559
rect 193 487 199 521
rect 233 487 239 521
rect 193 449 239 487
rect 193 415 199 449
rect 233 415 239 449
rect 193 377 239 415
rect 193 343 199 377
rect 233 343 239 377
rect 193 305 239 343
rect 193 271 199 305
rect 233 271 239 305
rect 193 233 239 271
rect 193 199 199 233
rect 233 199 239 233
rect 193 161 239 199
rect 193 127 199 161
rect 233 127 239 161
rect 193 89 239 127
rect 193 55 199 89
rect 233 55 239 89
rect 193 17 239 55
rect 193 -17 199 17
rect 233 -17 239 17
rect 193 -55 239 -17
rect 193 -89 199 -55
rect 233 -89 239 -55
rect 193 -127 239 -89
rect 193 -161 199 -127
rect 233 -161 239 -127
rect 193 -199 239 -161
rect 193 -233 199 -199
rect 233 -233 239 -199
rect 193 -271 239 -233
rect 193 -305 199 -271
rect 233 -305 239 -271
rect 193 -343 239 -305
rect 193 -377 199 -343
rect 233 -377 239 -343
rect 193 -415 239 -377
rect 193 -449 199 -415
rect 233 -449 239 -415
rect 193 -487 239 -449
rect 193 -521 199 -487
rect 233 -521 239 -487
rect 193 -559 239 -521
rect 193 -593 199 -559
rect 233 -593 239 -559
rect 193 -631 239 -593
rect 193 -665 199 -631
rect 233 -665 239 -631
rect 193 -703 239 -665
rect 193 -737 199 -703
rect 233 -737 239 -703
rect 193 -775 239 -737
rect 193 -809 199 -775
rect 233 -809 239 -775
rect 193 -847 239 -809
rect 193 -881 199 -847
rect 233 -881 239 -847
rect 193 -919 239 -881
rect 193 -953 199 -919
rect 233 -953 239 -919
rect 193 -991 239 -953
rect 193 -1025 199 -991
rect 233 -1025 239 -991
rect 193 -1063 239 -1025
rect 193 -1097 199 -1063
rect 233 -1097 239 -1063
rect 193 -1135 239 -1097
rect 193 -1169 199 -1135
rect 233 -1169 239 -1135
rect 193 -1207 239 -1169
rect 193 -1241 199 -1207
rect 233 -1241 239 -1207
rect 193 -1279 239 -1241
rect 193 -1313 199 -1279
rect 233 -1313 239 -1279
rect 193 -1351 239 -1313
rect 193 -1385 199 -1351
rect 233 -1385 239 -1351
rect 193 -1423 239 -1385
rect 193 -1457 199 -1423
rect 233 -1457 239 -1423
rect 193 -1495 239 -1457
rect 193 -1529 199 -1495
rect 233 -1529 239 -1495
rect 193 -1567 239 -1529
rect 193 -1601 199 -1567
rect 233 -1601 239 -1567
rect 193 -1639 239 -1601
rect 193 -1673 199 -1639
rect 233 -1673 239 -1639
rect 193 -1711 239 -1673
rect 193 -1745 199 -1711
rect 233 -1745 239 -1711
rect 193 -1783 239 -1745
rect 193 -1817 199 -1783
rect 233 -1817 239 -1783
rect 193 -1855 239 -1817
rect 193 -1889 199 -1855
rect 233 -1889 239 -1855
rect 193 -1927 239 -1889
rect 193 -1961 199 -1927
rect 233 -1961 239 -1927
rect 193 -1999 239 -1961
rect 193 -2033 199 -1999
rect 233 -2033 239 -1999
rect 193 -2071 239 -2033
rect 193 -2105 199 -2071
rect 233 -2105 239 -2071
rect 193 -2143 239 -2105
rect 193 -2177 199 -2143
rect 233 -2177 239 -2143
rect 193 -2215 239 -2177
rect 193 -2249 199 -2215
rect 233 -2249 239 -2215
rect 193 -2287 239 -2249
rect 193 -2321 199 -2287
rect 233 -2321 239 -2287
rect 193 -2359 239 -2321
rect 193 -2393 199 -2359
rect 233 -2393 239 -2359
rect 193 -2431 239 -2393
rect 193 -2465 199 -2431
rect 233 -2465 239 -2431
rect 193 -2500 239 -2465
rect 301 2465 347 2500
rect 301 2431 307 2465
rect 341 2431 347 2465
rect 301 2393 347 2431
rect 301 2359 307 2393
rect 341 2359 347 2393
rect 301 2321 347 2359
rect 301 2287 307 2321
rect 341 2287 347 2321
rect 301 2249 347 2287
rect 301 2215 307 2249
rect 341 2215 347 2249
rect 301 2177 347 2215
rect 301 2143 307 2177
rect 341 2143 347 2177
rect 301 2105 347 2143
rect 301 2071 307 2105
rect 341 2071 347 2105
rect 301 2033 347 2071
rect 301 1999 307 2033
rect 341 1999 347 2033
rect 301 1961 347 1999
rect 301 1927 307 1961
rect 341 1927 347 1961
rect 301 1889 347 1927
rect 301 1855 307 1889
rect 341 1855 347 1889
rect 301 1817 347 1855
rect 301 1783 307 1817
rect 341 1783 347 1817
rect 301 1745 347 1783
rect 301 1711 307 1745
rect 341 1711 347 1745
rect 301 1673 347 1711
rect 301 1639 307 1673
rect 341 1639 347 1673
rect 301 1601 347 1639
rect 301 1567 307 1601
rect 341 1567 347 1601
rect 301 1529 347 1567
rect 301 1495 307 1529
rect 341 1495 347 1529
rect 301 1457 347 1495
rect 301 1423 307 1457
rect 341 1423 347 1457
rect 301 1385 347 1423
rect 301 1351 307 1385
rect 341 1351 347 1385
rect 301 1313 347 1351
rect 301 1279 307 1313
rect 341 1279 347 1313
rect 301 1241 347 1279
rect 301 1207 307 1241
rect 341 1207 347 1241
rect 301 1169 347 1207
rect 301 1135 307 1169
rect 341 1135 347 1169
rect 301 1097 347 1135
rect 301 1063 307 1097
rect 341 1063 347 1097
rect 301 1025 347 1063
rect 301 991 307 1025
rect 341 991 347 1025
rect 301 953 347 991
rect 301 919 307 953
rect 341 919 347 953
rect 301 881 347 919
rect 301 847 307 881
rect 341 847 347 881
rect 301 809 347 847
rect 301 775 307 809
rect 341 775 347 809
rect 301 737 347 775
rect 301 703 307 737
rect 341 703 347 737
rect 301 665 347 703
rect 301 631 307 665
rect 341 631 347 665
rect 301 593 347 631
rect 301 559 307 593
rect 341 559 347 593
rect 301 521 347 559
rect 301 487 307 521
rect 341 487 347 521
rect 301 449 347 487
rect 301 415 307 449
rect 341 415 347 449
rect 301 377 347 415
rect 301 343 307 377
rect 341 343 347 377
rect 301 305 347 343
rect 301 271 307 305
rect 341 271 347 305
rect 301 233 347 271
rect 301 199 307 233
rect 341 199 347 233
rect 301 161 347 199
rect 301 127 307 161
rect 341 127 347 161
rect 301 89 347 127
rect 301 55 307 89
rect 341 55 347 89
rect 301 17 347 55
rect 301 -17 307 17
rect 341 -17 347 17
rect 301 -55 347 -17
rect 301 -89 307 -55
rect 341 -89 347 -55
rect 301 -127 347 -89
rect 301 -161 307 -127
rect 341 -161 347 -127
rect 301 -199 347 -161
rect 301 -233 307 -199
rect 341 -233 347 -199
rect 301 -271 347 -233
rect 301 -305 307 -271
rect 341 -305 347 -271
rect 301 -343 347 -305
rect 301 -377 307 -343
rect 341 -377 347 -343
rect 301 -415 347 -377
rect 301 -449 307 -415
rect 341 -449 347 -415
rect 301 -487 347 -449
rect 301 -521 307 -487
rect 341 -521 347 -487
rect 301 -559 347 -521
rect 301 -593 307 -559
rect 341 -593 347 -559
rect 301 -631 347 -593
rect 301 -665 307 -631
rect 341 -665 347 -631
rect 301 -703 347 -665
rect 301 -737 307 -703
rect 341 -737 347 -703
rect 301 -775 347 -737
rect 301 -809 307 -775
rect 341 -809 347 -775
rect 301 -847 347 -809
rect 301 -881 307 -847
rect 341 -881 347 -847
rect 301 -919 347 -881
rect 301 -953 307 -919
rect 341 -953 347 -919
rect 301 -991 347 -953
rect 301 -1025 307 -991
rect 341 -1025 347 -991
rect 301 -1063 347 -1025
rect 301 -1097 307 -1063
rect 341 -1097 347 -1063
rect 301 -1135 347 -1097
rect 301 -1169 307 -1135
rect 341 -1169 347 -1135
rect 301 -1207 347 -1169
rect 301 -1241 307 -1207
rect 341 -1241 347 -1207
rect 301 -1279 347 -1241
rect 301 -1313 307 -1279
rect 341 -1313 347 -1279
rect 301 -1351 347 -1313
rect 301 -1385 307 -1351
rect 341 -1385 347 -1351
rect 301 -1423 347 -1385
rect 301 -1457 307 -1423
rect 341 -1457 347 -1423
rect 301 -1495 347 -1457
rect 301 -1529 307 -1495
rect 341 -1529 347 -1495
rect 301 -1567 347 -1529
rect 301 -1601 307 -1567
rect 341 -1601 347 -1567
rect 301 -1639 347 -1601
rect 301 -1673 307 -1639
rect 341 -1673 347 -1639
rect 301 -1711 347 -1673
rect 301 -1745 307 -1711
rect 341 -1745 347 -1711
rect 301 -1783 347 -1745
rect 301 -1817 307 -1783
rect 341 -1817 347 -1783
rect 301 -1855 347 -1817
rect 301 -1889 307 -1855
rect 341 -1889 347 -1855
rect 301 -1927 347 -1889
rect 301 -1961 307 -1927
rect 341 -1961 347 -1927
rect 301 -1999 347 -1961
rect 301 -2033 307 -1999
rect 341 -2033 347 -1999
rect 301 -2071 347 -2033
rect 301 -2105 307 -2071
rect 341 -2105 347 -2071
rect 301 -2143 347 -2105
rect 301 -2177 307 -2143
rect 341 -2177 347 -2143
rect 301 -2215 347 -2177
rect 301 -2249 307 -2215
rect 341 -2249 347 -2215
rect 301 -2287 347 -2249
rect 301 -2321 307 -2287
rect 341 -2321 347 -2287
rect 301 -2359 347 -2321
rect 301 -2393 307 -2359
rect 341 -2393 347 -2359
rect 301 -2431 347 -2393
rect 301 -2465 307 -2431
rect 341 -2465 347 -2431
rect 301 -2500 347 -2465
rect 409 2465 455 2500
rect 409 2431 415 2465
rect 449 2431 455 2465
rect 409 2393 455 2431
rect 409 2359 415 2393
rect 449 2359 455 2393
rect 409 2321 455 2359
rect 409 2287 415 2321
rect 449 2287 455 2321
rect 409 2249 455 2287
rect 409 2215 415 2249
rect 449 2215 455 2249
rect 409 2177 455 2215
rect 409 2143 415 2177
rect 449 2143 455 2177
rect 409 2105 455 2143
rect 409 2071 415 2105
rect 449 2071 455 2105
rect 409 2033 455 2071
rect 409 1999 415 2033
rect 449 1999 455 2033
rect 409 1961 455 1999
rect 409 1927 415 1961
rect 449 1927 455 1961
rect 409 1889 455 1927
rect 409 1855 415 1889
rect 449 1855 455 1889
rect 409 1817 455 1855
rect 409 1783 415 1817
rect 449 1783 455 1817
rect 409 1745 455 1783
rect 409 1711 415 1745
rect 449 1711 455 1745
rect 409 1673 455 1711
rect 409 1639 415 1673
rect 449 1639 455 1673
rect 409 1601 455 1639
rect 409 1567 415 1601
rect 449 1567 455 1601
rect 409 1529 455 1567
rect 409 1495 415 1529
rect 449 1495 455 1529
rect 409 1457 455 1495
rect 409 1423 415 1457
rect 449 1423 455 1457
rect 409 1385 455 1423
rect 409 1351 415 1385
rect 449 1351 455 1385
rect 409 1313 455 1351
rect 409 1279 415 1313
rect 449 1279 455 1313
rect 409 1241 455 1279
rect 409 1207 415 1241
rect 449 1207 455 1241
rect 409 1169 455 1207
rect 409 1135 415 1169
rect 449 1135 455 1169
rect 409 1097 455 1135
rect 409 1063 415 1097
rect 449 1063 455 1097
rect 409 1025 455 1063
rect 409 991 415 1025
rect 449 991 455 1025
rect 409 953 455 991
rect 409 919 415 953
rect 449 919 455 953
rect 409 881 455 919
rect 409 847 415 881
rect 449 847 455 881
rect 409 809 455 847
rect 409 775 415 809
rect 449 775 455 809
rect 409 737 455 775
rect 409 703 415 737
rect 449 703 455 737
rect 409 665 455 703
rect 409 631 415 665
rect 449 631 455 665
rect 409 593 455 631
rect 409 559 415 593
rect 449 559 455 593
rect 409 521 455 559
rect 409 487 415 521
rect 449 487 455 521
rect 409 449 455 487
rect 409 415 415 449
rect 449 415 455 449
rect 409 377 455 415
rect 409 343 415 377
rect 449 343 455 377
rect 409 305 455 343
rect 409 271 415 305
rect 449 271 455 305
rect 409 233 455 271
rect 409 199 415 233
rect 449 199 455 233
rect 409 161 455 199
rect 409 127 415 161
rect 449 127 455 161
rect 409 89 455 127
rect 409 55 415 89
rect 449 55 455 89
rect 409 17 455 55
rect 409 -17 415 17
rect 449 -17 455 17
rect 409 -55 455 -17
rect 409 -89 415 -55
rect 449 -89 455 -55
rect 409 -127 455 -89
rect 409 -161 415 -127
rect 449 -161 455 -127
rect 409 -199 455 -161
rect 409 -233 415 -199
rect 449 -233 455 -199
rect 409 -271 455 -233
rect 409 -305 415 -271
rect 449 -305 455 -271
rect 409 -343 455 -305
rect 409 -377 415 -343
rect 449 -377 455 -343
rect 409 -415 455 -377
rect 409 -449 415 -415
rect 449 -449 455 -415
rect 409 -487 455 -449
rect 409 -521 415 -487
rect 449 -521 455 -487
rect 409 -559 455 -521
rect 409 -593 415 -559
rect 449 -593 455 -559
rect 409 -631 455 -593
rect 409 -665 415 -631
rect 449 -665 455 -631
rect 409 -703 455 -665
rect 409 -737 415 -703
rect 449 -737 455 -703
rect 409 -775 455 -737
rect 409 -809 415 -775
rect 449 -809 455 -775
rect 409 -847 455 -809
rect 409 -881 415 -847
rect 449 -881 455 -847
rect 409 -919 455 -881
rect 409 -953 415 -919
rect 449 -953 455 -919
rect 409 -991 455 -953
rect 409 -1025 415 -991
rect 449 -1025 455 -991
rect 409 -1063 455 -1025
rect 409 -1097 415 -1063
rect 449 -1097 455 -1063
rect 409 -1135 455 -1097
rect 409 -1169 415 -1135
rect 449 -1169 455 -1135
rect 409 -1207 455 -1169
rect 409 -1241 415 -1207
rect 449 -1241 455 -1207
rect 409 -1279 455 -1241
rect 409 -1313 415 -1279
rect 449 -1313 455 -1279
rect 409 -1351 455 -1313
rect 409 -1385 415 -1351
rect 449 -1385 455 -1351
rect 409 -1423 455 -1385
rect 409 -1457 415 -1423
rect 449 -1457 455 -1423
rect 409 -1495 455 -1457
rect 409 -1529 415 -1495
rect 449 -1529 455 -1495
rect 409 -1567 455 -1529
rect 409 -1601 415 -1567
rect 449 -1601 455 -1567
rect 409 -1639 455 -1601
rect 409 -1673 415 -1639
rect 449 -1673 455 -1639
rect 409 -1711 455 -1673
rect 409 -1745 415 -1711
rect 449 -1745 455 -1711
rect 409 -1783 455 -1745
rect 409 -1817 415 -1783
rect 449 -1817 455 -1783
rect 409 -1855 455 -1817
rect 409 -1889 415 -1855
rect 449 -1889 455 -1855
rect 409 -1927 455 -1889
rect 409 -1961 415 -1927
rect 449 -1961 455 -1927
rect 409 -1999 455 -1961
rect 409 -2033 415 -1999
rect 449 -2033 455 -1999
rect 409 -2071 455 -2033
rect 409 -2105 415 -2071
rect 449 -2105 455 -2071
rect 409 -2143 455 -2105
rect 409 -2177 415 -2143
rect 449 -2177 455 -2143
rect 409 -2215 455 -2177
rect 409 -2249 415 -2215
rect 449 -2249 455 -2215
rect 409 -2287 455 -2249
rect 409 -2321 415 -2287
rect 449 -2321 455 -2287
rect 409 -2359 455 -2321
rect 409 -2393 415 -2359
rect 449 -2393 455 -2359
rect 409 -2431 455 -2393
rect 409 -2465 415 -2431
rect 449 -2465 455 -2431
rect 409 -2500 455 -2465
rect -407 -2547 -349 -2541
rect -407 -2581 -395 -2547
rect -361 -2581 -349 -2547
rect -407 -2587 -349 -2581
rect -191 -2547 -133 -2541
rect -191 -2581 -179 -2547
rect -145 -2581 -133 -2547
rect -191 -2587 -133 -2581
rect 25 -2547 83 -2541
rect 25 -2581 37 -2547
rect 71 -2581 83 -2547
rect 25 -2587 83 -2581
rect 241 -2547 299 -2541
rect 241 -2581 253 -2547
rect 287 -2581 299 -2547
rect 241 -2587 299 -2581
<< properties >>
string FIXED_BBOX -546 -2666 546 2666
<< end >>
