** sch_path: /usr/local/share/pdk/sky130A/libs.tech/xschem/sky130_tests/test_ac.sch
**.subckt test_ac
XM1 G PLUS S GND sky130_fd_pr__nfet_01v8_lvt L=2 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 OUT MINUS S GND sky130_fd_pr__nfet_01v8_lvt L=2 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net3 BIAS GND GND sky130_fd_pr__nfet_01v8_lvt L=4 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 OUT G VCC VCC sky130_fd_pr__pfet_01v8_lvt L=4 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 G G VCC VCC sky130_fd_pr__pfet_01v8_lvt L=4 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vtail S net3 0
.save i(vtail)
V1 BIAS GND 0.7
V2 VCC GND 1.8
V3 PLUS GND 0.91
V4 IN GND 0 ac 1 0 sin(0 1m 100meg 0 0 0)
C2 MINUS IN 1T m=1
L1 OUT MINUS 1T m=1
E1 net1 GND S GND 1
XM6 net2 OUT net1 GND sky130_fd_pr__nfet_01v8_lvt L=2 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
E2 net2 GND OUT GND 1
**** begin user architecture code
.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt



.save
+ @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gm]
+ @m.xm2.msky130_fd_pr__nfet_01v8_lvt[gm]
+ @m.xm4.msky130_fd_pr__nfet_01v8_lvt[gm]
+ @m.xm3.msky130_fd_pr__pfet_01v8_lvt[gm]
+ @m.xm5.msky130_fd_pr__pfet_01v8_lvt[gm]
+ v(@m.xm5.msky130_fd_pr__pfet_01v8_lvt[vth])
+ @m.xm5.msky130_fd_pr__pfet_01v8_lvt[gds]
+ v(@m.xm3.msky130_fd_pr__pfet_01v8_lvt[vth])
+ @m.xm3.msky130_fd_pr__pfet_01v8_lvt[gds]

.option reltol=1e-5
+  abstol=1e-14 savecurrents
.control
  save all
  op
  remzerovec
  write test_ac.raw
  set appendwrite
  ac dec 10 1 1e12
  remzerovec
  write test_ac.raw
  tran 0.1n 100n
  write test_ac.raw
.endc






**** end user architecture code
**.ends
.end
