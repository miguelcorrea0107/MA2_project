** sch_path: /Users/miguelcorrea/Desktop/MA2_project/Amplifier_Inv/xschem/v2/tb_res.sch
**.subckt tb_res
VP VCC GND 1.125
Vin in out ac 1e-3 sin(0.8 0.001 5000 0 0 0)
Vdc out GND 0.53577
XM1 in VCC out GND sky130_fd_pr__nfet_01v8 L=20 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt



.control

  ac lin 100 1 100k
  save all
  let r = (v(out)-v(in))/i(Vin)
  write tb_inv_sky130_a_res_AC_v2.raw r

  tran 0.1u 4m
  save all
  write test.raw

  exit 0
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VCC
.end
