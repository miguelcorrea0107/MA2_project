** sch_path: /Users/miguelcorrea/Desktop/MA2_project/Amplifier_Inv/xschem/DC_tb.sch
**.subckt DC_tb
VN VSS GND 0
VP VCC GND 1.125
.save i(vp)
Vin in GND 0.44866 ac 1e-3 sin(0.44866 0.001 1000 0 0 0)
.save i(vin)
Rl out GND 1e60 m=1
x1 test in VCC VSS not W_N=250 L_N=1 W_P=180 L_P=0.25 m=1
XC2 out GND sky130_fd_pr__cap_mim_m3_1 W=50 L=50 MF=1 m=1
XR1 test in GND sky130_fd_pr__res_xhigh_po W=0.15 L=90000 mult=1 m=1
XR2 out test GND sky130_fd_pr__res_xhigh_po W=0.15 L=50 mult=1 m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt



.control

  dc Vin 0 1 0.00001
  save all v(in) v(out)
  write DC_tb.raw v(in) v(out)

.endc


**** end user architecture code
**.ends

* expanding   symbol:  sky130_tests/not.sym # of pins=2
** sym_path: /usr/local/share/pdk/sky130A/libs.tech/xschem/sky130_tests/not.sym
** sch_path: /usr/local/share/pdk/sky130A/libs.tech/xschem/sky130_tests/not.sch
.subckt not y a VCCPIN VSSPIN     W_N=1 L_N=0.15 W_P=2 L_P=0.15
*.opin y
*.ipin a
XM1 y a VSSPIN VSSPIN sky130_fd_pr__nfet_01v8 L=L_N W=W_N nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 y a VCCPIN VCCPIN sky130_fd_pr__pfet_01v8 L=L_P W=W_P nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.GLOBAL VSS
.GLOBAL VCC
.end
