** sch_path: /Users/miguelcorrea/Desktop/MA2_project/Amplifier_Inv/xschem/v2/tb_res.sch
**.subckt tb_res
Vgs gs net1 dc 1.125
Vds in net1 ac 1e-3
XM1 in gs net1 GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vs net1 GND dc 0.5
**** begin user architecture code

** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt



.control

  let start_vgs = 0.2
  let stop_vgs = 0.8
  let delta_vgs = 0.05
  let vgs_act = start_vgs

  while vgs_act le stop_vgs
  alter vgs dc vgs_act
  ac dec 100 0.1 100k
  let r = v(in)/(-i(Vds))
  save all
  write tb_inv_sky130_a_res_AC_v2.raw r
  set appendwrite
  let vgs_act = vgs_act + delta_vgs
  end

.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
