** sch_path: /Users/miguelcorrea/Desktop/MA2_project/Amplifier_Inv/xschem/v4/tb_inv_sky130_a_v4.sch
**.subckt tb_inv_sky130_a_v4
VN VSS GND 0
VP VCC GND dc 1.125
.save i(vp)
Vin in GND 0.48731 ac 1e-3 sin(0.48731 0.001 5000 0 0 0)
.save i(vin)
Rl out GND 1e60 m=1
VG2 net1 GND dc 1.085
VG1 net2 GND dc 0.725
x1 net2 VCC net1 out in VSS inv_sky130_a_v4
**** begin user architecture code

** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt



.control

  op
  save all
  let gmn = @m.x1.xm4.msky130_fd_pr__nfet_01v8[gm]
  let gmp = @m.x1.xm5'.msky130_fd_pr__pfet_01v8[gm]
  let gdsn = @m.x1.xm4.msky130_fd_pr__nfet_01v8[gds]
  let gdsp = @m.x1.xm5.msky130_fd_pr__pfet_01v8[gds]
  let cgsn = @m.x1.xm4.msky130_fd_pr__nfet_01v8[cgs]
  let cgsp = @m.x1.xm5.msky130_fd_pr__pfet_01v8[cgs]
  let cgdn = @m.x1.xm4.msky130_fd_pr__nfet_01v8[cgd]
  let cgdp = @m.x1.xm5.msky130_fd_pr__pfet_01v8[cgd]
  write tb_inv_sky130_a_op_v4.raw gmn gmp gdsn gdsp cgsn cgsp cgdn cgdp

  ac dec 1000 1 1e8
  save all
  let gain = db(v(out)/v(in))
  let gain_vs1 = db(v(x1.vs1)/v(in))
  let phase = phase(v(out)/v(in))
  write tb_inv_sky130_a_AC_v4.raw gain gain_vs1

  noise v(out) Vin dec 1000 300 10k 10
  save all
  write tb_inv_sky130_a_noise_v4.raw

  noise v(out) Vin dec 1000 300 10k
  save all
  setplot noise1
  write tb_inv_sky130_a_noise_spectrum_v4.raw

  dc Vin 0 1.125 0.00001
  save all v(out) v(x1.vs1) v(x1.vd1)
  write tb_inv_sky130_a_DC_v4.raw v(out) v(x1.vs1) v(x1.vd1)

  tran 0.1u 4m
  save all
  let pw_in = i(Vin)*v(in)
  let pw_vcc = i(Vp)*1.125
  let pw_vg1 = i(Vg1)*0.725
  let pw_vg2 = i(Vg2)*1.085
  let pw_total = pw_in+pw_vcc
  meas tran avg_pw_total AVG pw_total FROM=0 TO=2m
  meas tran avg_pw_in AVG pw_in FROM=0 TO=2m
  meas tran avg_pw_vcc AVG pw_vcc FROM=0 TO=2m
  write tb_inv_sky130_a_tran_v4.raw v(in) v(out) v(x1.vd1) v(x1.vs1) v(vg1) v(vg2) avg_pw_total

  exit 0
.endc


**** end user architecture code
**.ends

* expanding   symbol:  v4/inv_sky130_a_v4.sym # of pins=6
** sym_path: /Users/miguelcorrea/Desktop/MA2_project/Amplifier_Inv/xschem/v4/inv_sky130_a_v4.sym
** sch_path: /Users/miguelcorrea/Desktop/MA2_project/Amplifier_Inv/xschem/v4/inv_sky130_a_v4.sch
.subckt inv_sky130_a_v4 VG1 VCC VG2 out in VSS
*.ipin in
*.opin out
*.ipin VG1
*.ipin VG2
*.ipin VSS
*.ipin VCC
XC1 in VD1 sky130_fd_pr__cap_mim_m3_1 W=26 L=26 MF=1 m=1
XM1 VD1 VG1 VS1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)
+ * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 VS1 VG2 out VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)
+ * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 VSS out VSS VSS sky130_fd_pr__nfet_01v8 L=10 W=100 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)
+ * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 VS1 VD1 VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=250 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)
+ * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 VS1 VD1 VCC VCC sky130_fd_pr__pfet_01v8 L=0.25 W=200 nf=8 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)
+ * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
