magic
tech sky130A
magscale 1 2
timestamp 1716644424
<< pwell >>
rect -4273 -2700 4273 2700
<< nmos >>
rect -4087 -2500 -2087 2500
rect -2029 -2500 -29 2500
rect 29 -2500 2029 2500
rect 2087 -2500 4087 2500
<< ndiff >>
rect -4145 2465 -4087 2500
rect -4145 2431 -4133 2465
rect -4099 2431 -4087 2465
rect -4145 2397 -4087 2431
rect -4145 2363 -4133 2397
rect -4099 2363 -4087 2397
rect -4145 2329 -4087 2363
rect -4145 2295 -4133 2329
rect -4099 2295 -4087 2329
rect -4145 2261 -4087 2295
rect -4145 2227 -4133 2261
rect -4099 2227 -4087 2261
rect -4145 2193 -4087 2227
rect -4145 2159 -4133 2193
rect -4099 2159 -4087 2193
rect -4145 2125 -4087 2159
rect -4145 2091 -4133 2125
rect -4099 2091 -4087 2125
rect -4145 2057 -4087 2091
rect -4145 2023 -4133 2057
rect -4099 2023 -4087 2057
rect -4145 1989 -4087 2023
rect -4145 1955 -4133 1989
rect -4099 1955 -4087 1989
rect -4145 1921 -4087 1955
rect -4145 1887 -4133 1921
rect -4099 1887 -4087 1921
rect -4145 1853 -4087 1887
rect -4145 1819 -4133 1853
rect -4099 1819 -4087 1853
rect -4145 1785 -4087 1819
rect -4145 1751 -4133 1785
rect -4099 1751 -4087 1785
rect -4145 1717 -4087 1751
rect -4145 1683 -4133 1717
rect -4099 1683 -4087 1717
rect -4145 1649 -4087 1683
rect -4145 1615 -4133 1649
rect -4099 1615 -4087 1649
rect -4145 1581 -4087 1615
rect -4145 1547 -4133 1581
rect -4099 1547 -4087 1581
rect -4145 1513 -4087 1547
rect -4145 1479 -4133 1513
rect -4099 1479 -4087 1513
rect -4145 1445 -4087 1479
rect -4145 1411 -4133 1445
rect -4099 1411 -4087 1445
rect -4145 1377 -4087 1411
rect -4145 1343 -4133 1377
rect -4099 1343 -4087 1377
rect -4145 1309 -4087 1343
rect -4145 1275 -4133 1309
rect -4099 1275 -4087 1309
rect -4145 1241 -4087 1275
rect -4145 1207 -4133 1241
rect -4099 1207 -4087 1241
rect -4145 1173 -4087 1207
rect -4145 1139 -4133 1173
rect -4099 1139 -4087 1173
rect -4145 1105 -4087 1139
rect -4145 1071 -4133 1105
rect -4099 1071 -4087 1105
rect -4145 1037 -4087 1071
rect -4145 1003 -4133 1037
rect -4099 1003 -4087 1037
rect -4145 969 -4087 1003
rect -4145 935 -4133 969
rect -4099 935 -4087 969
rect -4145 901 -4087 935
rect -4145 867 -4133 901
rect -4099 867 -4087 901
rect -4145 833 -4087 867
rect -4145 799 -4133 833
rect -4099 799 -4087 833
rect -4145 765 -4087 799
rect -4145 731 -4133 765
rect -4099 731 -4087 765
rect -4145 697 -4087 731
rect -4145 663 -4133 697
rect -4099 663 -4087 697
rect -4145 629 -4087 663
rect -4145 595 -4133 629
rect -4099 595 -4087 629
rect -4145 561 -4087 595
rect -4145 527 -4133 561
rect -4099 527 -4087 561
rect -4145 493 -4087 527
rect -4145 459 -4133 493
rect -4099 459 -4087 493
rect -4145 425 -4087 459
rect -4145 391 -4133 425
rect -4099 391 -4087 425
rect -4145 357 -4087 391
rect -4145 323 -4133 357
rect -4099 323 -4087 357
rect -4145 289 -4087 323
rect -4145 255 -4133 289
rect -4099 255 -4087 289
rect -4145 221 -4087 255
rect -4145 187 -4133 221
rect -4099 187 -4087 221
rect -4145 153 -4087 187
rect -4145 119 -4133 153
rect -4099 119 -4087 153
rect -4145 85 -4087 119
rect -4145 51 -4133 85
rect -4099 51 -4087 85
rect -4145 17 -4087 51
rect -4145 -17 -4133 17
rect -4099 -17 -4087 17
rect -4145 -51 -4087 -17
rect -4145 -85 -4133 -51
rect -4099 -85 -4087 -51
rect -4145 -119 -4087 -85
rect -4145 -153 -4133 -119
rect -4099 -153 -4087 -119
rect -4145 -187 -4087 -153
rect -4145 -221 -4133 -187
rect -4099 -221 -4087 -187
rect -4145 -255 -4087 -221
rect -4145 -289 -4133 -255
rect -4099 -289 -4087 -255
rect -4145 -323 -4087 -289
rect -4145 -357 -4133 -323
rect -4099 -357 -4087 -323
rect -4145 -391 -4087 -357
rect -4145 -425 -4133 -391
rect -4099 -425 -4087 -391
rect -4145 -459 -4087 -425
rect -4145 -493 -4133 -459
rect -4099 -493 -4087 -459
rect -4145 -527 -4087 -493
rect -4145 -561 -4133 -527
rect -4099 -561 -4087 -527
rect -4145 -595 -4087 -561
rect -4145 -629 -4133 -595
rect -4099 -629 -4087 -595
rect -4145 -663 -4087 -629
rect -4145 -697 -4133 -663
rect -4099 -697 -4087 -663
rect -4145 -731 -4087 -697
rect -4145 -765 -4133 -731
rect -4099 -765 -4087 -731
rect -4145 -799 -4087 -765
rect -4145 -833 -4133 -799
rect -4099 -833 -4087 -799
rect -4145 -867 -4087 -833
rect -4145 -901 -4133 -867
rect -4099 -901 -4087 -867
rect -4145 -935 -4087 -901
rect -4145 -969 -4133 -935
rect -4099 -969 -4087 -935
rect -4145 -1003 -4087 -969
rect -4145 -1037 -4133 -1003
rect -4099 -1037 -4087 -1003
rect -4145 -1071 -4087 -1037
rect -4145 -1105 -4133 -1071
rect -4099 -1105 -4087 -1071
rect -4145 -1139 -4087 -1105
rect -4145 -1173 -4133 -1139
rect -4099 -1173 -4087 -1139
rect -4145 -1207 -4087 -1173
rect -4145 -1241 -4133 -1207
rect -4099 -1241 -4087 -1207
rect -4145 -1275 -4087 -1241
rect -4145 -1309 -4133 -1275
rect -4099 -1309 -4087 -1275
rect -4145 -1343 -4087 -1309
rect -4145 -1377 -4133 -1343
rect -4099 -1377 -4087 -1343
rect -4145 -1411 -4087 -1377
rect -4145 -1445 -4133 -1411
rect -4099 -1445 -4087 -1411
rect -4145 -1479 -4087 -1445
rect -4145 -1513 -4133 -1479
rect -4099 -1513 -4087 -1479
rect -4145 -1547 -4087 -1513
rect -4145 -1581 -4133 -1547
rect -4099 -1581 -4087 -1547
rect -4145 -1615 -4087 -1581
rect -4145 -1649 -4133 -1615
rect -4099 -1649 -4087 -1615
rect -4145 -1683 -4087 -1649
rect -4145 -1717 -4133 -1683
rect -4099 -1717 -4087 -1683
rect -4145 -1751 -4087 -1717
rect -4145 -1785 -4133 -1751
rect -4099 -1785 -4087 -1751
rect -4145 -1819 -4087 -1785
rect -4145 -1853 -4133 -1819
rect -4099 -1853 -4087 -1819
rect -4145 -1887 -4087 -1853
rect -4145 -1921 -4133 -1887
rect -4099 -1921 -4087 -1887
rect -4145 -1955 -4087 -1921
rect -4145 -1989 -4133 -1955
rect -4099 -1989 -4087 -1955
rect -4145 -2023 -4087 -1989
rect -4145 -2057 -4133 -2023
rect -4099 -2057 -4087 -2023
rect -4145 -2091 -4087 -2057
rect -4145 -2125 -4133 -2091
rect -4099 -2125 -4087 -2091
rect -4145 -2159 -4087 -2125
rect -4145 -2193 -4133 -2159
rect -4099 -2193 -4087 -2159
rect -4145 -2227 -4087 -2193
rect -4145 -2261 -4133 -2227
rect -4099 -2261 -4087 -2227
rect -4145 -2295 -4087 -2261
rect -4145 -2329 -4133 -2295
rect -4099 -2329 -4087 -2295
rect -4145 -2363 -4087 -2329
rect -4145 -2397 -4133 -2363
rect -4099 -2397 -4087 -2363
rect -4145 -2431 -4087 -2397
rect -4145 -2465 -4133 -2431
rect -4099 -2465 -4087 -2431
rect -4145 -2500 -4087 -2465
rect -2087 2465 -2029 2500
rect -2087 2431 -2075 2465
rect -2041 2431 -2029 2465
rect -2087 2397 -2029 2431
rect -2087 2363 -2075 2397
rect -2041 2363 -2029 2397
rect -2087 2329 -2029 2363
rect -2087 2295 -2075 2329
rect -2041 2295 -2029 2329
rect -2087 2261 -2029 2295
rect -2087 2227 -2075 2261
rect -2041 2227 -2029 2261
rect -2087 2193 -2029 2227
rect -2087 2159 -2075 2193
rect -2041 2159 -2029 2193
rect -2087 2125 -2029 2159
rect -2087 2091 -2075 2125
rect -2041 2091 -2029 2125
rect -2087 2057 -2029 2091
rect -2087 2023 -2075 2057
rect -2041 2023 -2029 2057
rect -2087 1989 -2029 2023
rect -2087 1955 -2075 1989
rect -2041 1955 -2029 1989
rect -2087 1921 -2029 1955
rect -2087 1887 -2075 1921
rect -2041 1887 -2029 1921
rect -2087 1853 -2029 1887
rect -2087 1819 -2075 1853
rect -2041 1819 -2029 1853
rect -2087 1785 -2029 1819
rect -2087 1751 -2075 1785
rect -2041 1751 -2029 1785
rect -2087 1717 -2029 1751
rect -2087 1683 -2075 1717
rect -2041 1683 -2029 1717
rect -2087 1649 -2029 1683
rect -2087 1615 -2075 1649
rect -2041 1615 -2029 1649
rect -2087 1581 -2029 1615
rect -2087 1547 -2075 1581
rect -2041 1547 -2029 1581
rect -2087 1513 -2029 1547
rect -2087 1479 -2075 1513
rect -2041 1479 -2029 1513
rect -2087 1445 -2029 1479
rect -2087 1411 -2075 1445
rect -2041 1411 -2029 1445
rect -2087 1377 -2029 1411
rect -2087 1343 -2075 1377
rect -2041 1343 -2029 1377
rect -2087 1309 -2029 1343
rect -2087 1275 -2075 1309
rect -2041 1275 -2029 1309
rect -2087 1241 -2029 1275
rect -2087 1207 -2075 1241
rect -2041 1207 -2029 1241
rect -2087 1173 -2029 1207
rect -2087 1139 -2075 1173
rect -2041 1139 -2029 1173
rect -2087 1105 -2029 1139
rect -2087 1071 -2075 1105
rect -2041 1071 -2029 1105
rect -2087 1037 -2029 1071
rect -2087 1003 -2075 1037
rect -2041 1003 -2029 1037
rect -2087 969 -2029 1003
rect -2087 935 -2075 969
rect -2041 935 -2029 969
rect -2087 901 -2029 935
rect -2087 867 -2075 901
rect -2041 867 -2029 901
rect -2087 833 -2029 867
rect -2087 799 -2075 833
rect -2041 799 -2029 833
rect -2087 765 -2029 799
rect -2087 731 -2075 765
rect -2041 731 -2029 765
rect -2087 697 -2029 731
rect -2087 663 -2075 697
rect -2041 663 -2029 697
rect -2087 629 -2029 663
rect -2087 595 -2075 629
rect -2041 595 -2029 629
rect -2087 561 -2029 595
rect -2087 527 -2075 561
rect -2041 527 -2029 561
rect -2087 493 -2029 527
rect -2087 459 -2075 493
rect -2041 459 -2029 493
rect -2087 425 -2029 459
rect -2087 391 -2075 425
rect -2041 391 -2029 425
rect -2087 357 -2029 391
rect -2087 323 -2075 357
rect -2041 323 -2029 357
rect -2087 289 -2029 323
rect -2087 255 -2075 289
rect -2041 255 -2029 289
rect -2087 221 -2029 255
rect -2087 187 -2075 221
rect -2041 187 -2029 221
rect -2087 153 -2029 187
rect -2087 119 -2075 153
rect -2041 119 -2029 153
rect -2087 85 -2029 119
rect -2087 51 -2075 85
rect -2041 51 -2029 85
rect -2087 17 -2029 51
rect -2087 -17 -2075 17
rect -2041 -17 -2029 17
rect -2087 -51 -2029 -17
rect -2087 -85 -2075 -51
rect -2041 -85 -2029 -51
rect -2087 -119 -2029 -85
rect -2087 -153 -2075 -119
rect -2041 -153 -2029 -119
rect -2087 -187 -2029 -153
rect -2087 -221 -2075 -187
rect -2041 -221 -2029 -187
rect -2087 -255 -2029 -221
rect -2087 -289 -2075 -255
rect -2041 -289 -2029 -255
rect -2087 -323 -2029 -289
rect -2087 -357 -2075 -323
rect -2041 -357 -2029 -323
rect -2087 -391 -2029 -357
rect -2087 -425 -2075 -391
rect -2041 -425 -2029 -391
rect -2087 -459 -2029 -425
rect -2087 -493 -2075 -459
rect -2041 -493 -2029 -459
rect -2087 -527 -2029 -493
rect -2087 -561 -2075 -527
rect -2041 -561 -2029 -527
rect -2087 -595 -2029 -561
rect -2087 -629 -2075 -595
rect -2041 -629 -2029 -595
rect -2087 -663 -2029 -629
rect -2087 -697 -2075 -663
rect -2041 -697 -2029 -663
rect -2087 -731 -2029 -697
rect -2087 -765 -2075 -731
rect -2041 -765 -2029 -731
rect -2087 -799 -2029 -765
rect -2087 -833 -2075 -799
rect -2041 -833 -2029 -799
rect -2087 -867 -2029 -833
rect -2087 -901 -2075 -867
rect -2041 -901 -2029 -867
rect -2087 -935 -2029 -901
rect -2087 -969 -2075 -935
rect -2041 -969 -2029 -935
rect -2087 -1003 -2029 -969
rect -2087 -1037 -2075 -1003
rect -2041 -1037 -2029 -1003
rect -2087 -1071 -2029 -1037
rect -2087 -1105 -2075 -1071
rect -2041 -1105 -2029 -1071
rect -2087 -1139 -2029 -1105
rect -2087 -1173 -2075 -1139
rect -2041 -1173 -2029 -1139
rect -2087 -1207 -2029 -1173
rect -2087 -1241 -2075 -1207
rect -2041 -1241 -2029 -1207
rect -2087 -1275 -2029 -1241
rect -2087 -1309 -2075 -1275
rect -2041 -1309 -2029 -1275
rect -2087 -1343 -2029 -1309
rect -2087 -1377 -2075 -1343
rect -2041 -1377 -2029 -1343
rect -2087 -1411 -2029 -1377
rect -2087 -1445 -2075 -1411
rect -2041 -1445 -2029 -1411
rect -2087 -1479 -2029 -1445
rect -2087 -1513 -2075 -1479
rect -2041 -1513 -2029 -1479
rect -2087 -1547 -2029 -1513
rect -2087 -1581 -2075 -1547
rect -2041 -1581 -2029 -1547
rect -2087 -1615 -2029 -1581
rect -2087 -1649 -2075 -1615
rect -2041 -1649 -2029 -1615
rect -2087 -1683 -2029 -1649
rect -2087 -1717 -2075 -1683
rect -2041 -1717 -2029 -1683
rect -2087 -1751 -2029 -1717
rect -2087 -1785 -2075 -1751
rect -2041 -1785 -2029 -1751
rect -2087 -1819 -2029 -1785
rect -2087 -1853 -2075 -1819
rect -2041 -1853 -2029 -1819
rect -2087 -1887 -2029 -1853
rect -2087 -1921 -2075 -1887
rect -2041 -1921 -2029 -1887
rect -2087 -1955 -2029 -1921
rect -2087 -1989 -2075 -1955
rect -2041 -1989 -2029 -1955
rect -2087 -2023 -2029 -1989
rect -2087 -2057 -2075 -2023
rect -2041 -2057 -2029 -2023
rect -2087 -2091 -2029 -2057
rect -2087 -2125 -2075 -2091
rect -2041 -2125 -2029 -2091
rect -2087 -2159 -2029 -2125
rect -2087 -2193 -2075 -2159
rect -2041 -2193 -2029 -2159
rect -2087 -2227 -2029 -2193
rect -2087 -2261 -2075 -2227
rect -2041 -2261 -2029 -2227
rect -2087 -2295 -2029 -2261
rect -2087 -2329 -2075 -2295
rect -2041 -2329 -2029 -2295
rect -2087 -2363 -2029 -2329
rect -2087 -2397 -2075 -2363
rect -2041 -2397 -2029 -2363
rect -2087 -2431 -2029 -2397
rect -2087 -2465 -2075 -2431
rect -2041 -2465 -2029 -2431
rect -2087 -2500 -2029 -2465
rect -29 2465 29 2500
rect -29 2431 -17 2465
rect 17 2431 29 2465
rect -29 2397 29 2431
rect -29 2363 -17 2397
rect 17 2363 29 2397
rect -29 2329 29 2363
rect -29 2295 -17 2329
rect 17 2295 29 2329
rect -29 2261 29 2295
rect -29 2227 -17 2261
rect 17 2227 29 2261
rect -29 2193 29 2227
rect -29 2159 -17 2193
rect 17 2159 29 2193
rect -29 2125 29 2159
rect -29 2091 -17 2125
rect 17 2091 29 2125
rect -29 2057 29 2091
rect -29 2023 -17 2057
rect 17 2023 29 2057
rect -29 1989 29 2023
rect -29 1955 -17 1989
rect 17 1955 29 1989
rect -29 1921 29 1955
rect -29 1887 -17 1921
rect 17 1887 29 1921
rect -29 1853 29 1887
rect -29 1819 -17 1853
rect 17 1819 29 1853
rect -29 1785 29 1819
rect -29 1751 -17 1785
rect 17 1751 29 1785
rect -29 1717 29 1751
rect -29 1683 -17 1717
rect 17 1683 29 1717
rect -29 1649 29 1683
rect -29 1615 -17 1649
rect 17 1615 29 1649
rect -29 1581 29 1615
rect -29 1547 -17 1581
rect 17 1547 29 1581
rect -29 1513 29 1547
rect -29 1479 -17 1513
rect 17 1479 29 1513
rect -29 1445 29 1479
rect -29 1411 -17 1445
rect 17 1411 29 1445
rect -29 1377 29 1411
rect -29 1343 -17 1377
rect 17 1343 29 1377
rect -29 1309 29 1343
rect -29 1275 -17 1309
rect 17 1275 29 1309
rect -29 1241 29 1275
rect -29 1207 -17 1241
rect 17 1207 29 1241
rect -29 1173 29 1207
rect -29 1139 -17 1173
rect 17 1139 29 1173
rect -29 1105 29 1139
rect -29 1071 -17 1105
rect 17 1071 29 1105
rect -29 1037 29 1071
rect -29 1003 -17 1037
rect 17 1003 29 1037
rect -29 969 29 1003
rect -29 935 -17 969
rect 17 935 29 969
rect -29 901 29 935
rect -29 867 -17 901
rect 17 867 29 901
rect -29 833 29 867
rect -29 799 -17 833
rect 17 799 29 833
rect -29 765 29 799
rect -29 731 -17 765
rect 17 731 29 765
rect -29 697 29 731
rect -29 663 -17 697
rect 17 663 29 697
rect -29 629 29 663
rect -29 595 -17 629
rect 17 595 29 629
rect -29 561 29 595
rect -29 527 -17 561
rect 17 527 29 561
rect -29 493 29 527
rect -29 459 -17 493
rect 17 459 29 493
rect -29 425 29 459
rect -29 391 -17 425
rect 17 391 29 425
rect -29 357 29 391
rect -29 323 -17 357
rect 17 323 29 357
rect -29 289 29 323
rect -29 255 -17 289
rect 17 255 29 289
rect -29 221 29 255
rect -29 187 -17 221
rect 17 187 29 221
rect -29 153 29 187
rect -29 119 -17 153
rect 17 119 29 153
rect -29 85 29 119
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -119 29 -85
rect -29 -153 -17 -119
rect 17 -153 29 -119
rect -29 -187 29 -153
rect -29 -221 -17 -187
rect 17 -221 29 -187
rect -29 -255 29 -221
rect -29 -289 -17 -255
rect 17 -289 29 -255
rect -29 -323 29 -289
rect -29 -357 -17 -323
rect 17 -357 29 -323
rect -29 -391 29 -357
rect -29 -425 -17 -391
rect 17 -425 29 -391
rect -29 -459 29 -425
rect -29 -493 -17 -459
rect 17 -493 29 -459
rect -29 -527 29 -493
rect -29 -561 -17 -527
rect 17 -561 29 -527
rect -29 -595 29 -561
rect -29 -629 -17 -595
rect 17 -629 29 -595
rect -29 -663 29 -629
rect -29 -697 -17 -663
rect 17 -697 29 -663
rect -29 -731 29 -697
rect -29 -765 -17 -731
rect 17 -765 29 -731
rect -29 -799 29 -765
rect -29 -833 -17 -799
rect 17 -833 29 -799
rect -29 -867 29 -833
rect -29 -901 -17 -867
rect 17 -901 29 -867
rect -29 -935 29 -901
rect -29 -969 -17 -935
rect 17 -969 29 -935
rect -29 -1003 29 -969
rect -29 -1037 -17 -1003
rect 17 -1037 29 -1003
rect -29 -1071 29 -1037
rect -29 -1105 -17 -1071
rect 17 -1105 29 -1071
rect -29 -1139 29 -1105
rect -29 -1173 -17 -1139
rect 17 -1173 29 -1139
rect -29 -1207 29 -1173
rect -29 -1241 -17 -1207
rect 17 -1241 29 -1207
rect -29 -1275 29 -1241
rect -29 -1309 -17 -1275
rect 17 -1309 29 -1275
rect -29 -1343 29 -1309
rect -29 -1377 -17 -1343
rect 17 -1377 29 -1343
rect -29 -1411 29 -1377
rect -29 -1445 -17 -1411
rect 17 -1445 29 -1411
rect -29 -1479 29 -1445
rect -29 -1513 -17 -1479
rect 17 -1513 29 -1479
rect -29 -1547 29 -1513
rect -29 -1581 -17 -1547
rect 17 -1581 29 -1547
rect -29 -1615 29 -1581
rect -29 -1649 -17 -1615
rect 17 -1649 29 -1615
rect -29 -1683 29 -1649
rect -29 -1717 -17 -1683
rect 17 -1717 29 -1683
rect -29 -1751 29 -1717
rect -29 -1785 -17 -1751
rect 17 -1785 29 -1751
rect -29 -1819 29 -1785
rect -29 -1853 -17 -1819
rect 17 -1853 29 -1819
rect -29 -1887 29 -1853
rect -29 -1921 -17 -1887
rect 17 -1921 29 -1887
rect -29 -1955 29 -1921
rect -29 -1989 -17 -1955
rect 17 -1989 29 -1955
rect -29 -2023 29 -1989
rect -29 -2057 -17 -2023
rect 17 -2057 29 -2023
rect -29 -2091 29 -2057
rect -29 -2125 -17 -2091
rect 17 -2125 29 -2091
rect -29 -2159 29 -2125
rect -29 -2193 -17 -2159
rect 17 -2193 29 -2159
rect -29 -2227 29 -2193
rect -29 -2261 -17 -2227
rect 17 -2261 29 -2227
rect -29 -2295 29 -2261
rect -29 -2329 -17 -2295
rect 17 -2329 29 -2295
rect -29 -2363 29 -2329
rect -29 -2397 -17 -2363
rect 17 -2397 29 -2363
rect -29 -2431 29 -2397
rect -29 -2465 -17 -2431
rect 17 -2465 29 -2431
rect -29 -2500 29 -2465
rect 2029 2465 2087 2500
rect 2029 2431 2041 2465
rect 2075 2431 2087 2465
rect 2029 2397 2087 2431
rect 2029 2363 2041 2397
rect 2075 2363 2087 2397
rect 2029 2329 2087 2363
rect 2029 2295 2041 2329
rect 2075 2295 2087 2329
rect 2029 2261 2087 2295
rect 2029 2227 2041 2261
rect 2075 2227 2087 2261
rect 2029 2193 2087 2227
rect 2029 2159 2041 2193
rect 2075 2159 2087 2193
rect 2029 2125 2087 2159
rect 2029 2091 2041 2125
rect 2075 2091 2087 2125
rect 2029 2057 2087 2091
rect 2029 2023 2041 2057
rect 2075 2023 2087 2057
rect 2029 1989 2087 2023
rect 2029 1955 2041 1989
rect 2075 1955 2087 1989
rect 2029 1921 2087 1955
rect 2029 1887 2041 1921
rect 2075 1887 2087 1921
rect 2029 1853 2087 1887
rect 2029 1819 2041 1853
rect 2075 1819 2087 1853
rect 2029 1785 2087 1819
rect 2029 1751 2041 1785
rect 2075 1751 2087 1785
rect 2029 1717 2087 1751
rect 2029 1683 2041 1717
rect 2075 1683 2087 1717
rect 2029 1649 2087 1683
rect 2029 1615 2041 1649
rect 2075 1615 2087 1649
rect 2029 1581 2087 1615
rect 2029 1547 2041 1581
rect 2075 1547 2087 1581
rect 2029 1513 2087 1547
rect 2029 1479 2041 1513
rect 2075 1479 2087 1513
rect 2029 1445 2087 1479
rect 2029 1411 2041 1445
rect 2075 1411 2087 1445
rect 2029 1377 2087 1411
rect 2029 1343 2041 1377
rect 2075 1343 2087 1377
rect 2029 1309 2087 1343
rect 2029 1275 2041 1309
rect 2075 1275 2087 1309
rect 2029 1241 2087 1275
rect 2029 1207 2041 1241
rect 2075 1207 2087 1241
rect 2029 1173 2087 1207
rect 2029 1139 2041 1173
rect 2075 1139 2087 1173
rect 2029 1105 2087 1139
rect 2029 1071 2041 1105
rect 2075 1071 2087 1105
rect 2029 1037 2087 1071
rect 2029 1003 2041 1037
rect 2075 1003 2087 1037
rect 2029 969 2087 1003
rect 2029 935 2041 969
rect 2075 935 2087 969
rect 2029 901 2087 935
rect 2029 867 2041 901
rect 2075 867 2087 901
rect 2029 833 2087 867
rect 2029 799 2041 833
rect 2075 799 2087 833
rect 2029 765 2087 799
rect 2029 731 2041 765
rect 2075 731 2087 765
rect 2029 697 2087 731
rect 2029 663 2041 697
rect 2075 663 2087 697
rect 2029 629 2087 663
rect 2029 595 2041 629
rect 2075 595 2087 629
rect 2029 561 2087 595
rect 2029 527 2041 561
rect 2075 527 2087 561
rect 2029 493 2087 527
rect 2029 459 2041 493
rect 2075 459 2087 493
rect 2029 425 2087 459
rect 2029 391 2041 425
rect 2075 391 2087 425
rect 2029 357 2087 391
rect 2029 323 2041 357
rect 2075 323 2087 357
rect 2029 289 2087 323
rect 2029 255 2041 289
rect 2075 255 2087 289
rect 2029 221 2087 255
rect 2029 187 2041 221
rect 2075 187 2087 221
rect 2029 153 2087 187
rect 2029 119 2041 153
rect 2075 119 2087 153
rect 2029 85 2087 119
rect 2029 51 2041 85
rect 2075 51 2087 85
rect 2029 17 2087 51
rect 2029 -17 2041 17
rect 2075 -17 2087 17
rect 2029 -51 2087 -17
rect 2029 -85 2041 -51
rect 2075 -85 2087 -51
rect 2029 -119 2087 -85
rect 2029 -153 2041 -119
rect 2075 -153 2087 -119
rect 2029 -187 2087 -153
rect 2029 -221 2041 -187
rect 2075 -221 2087 -187
rect 2029 -255 2087 -221
rect 2029 -289 2041 -255
rect 2075 -289 2087 -255
rect 2029 -323 2087 -289
rect 2029 -357 2041 -323
rect 2075 -357 2087 -323
rect 2029 -391 2087 -357
rect 2029 -425 2041 -391
rect 2075 -425 2087 -391
rect 2029 -459 2087 -425
rect 2029 -493 2041 -459
rect 2075 -493 2087 -459
rect 2029 -527 2087 -493
rect 2029 -561 2041 -527
rect 2075 -561 2087 -527
rect 2029 -595 2087 -561
rect 2029 -629 2041 -595
rect 2075 -629 2087 -595
rect 2029 -663 2087 -629
rect 2029 -697 2041 -663
rect 2075 -697 2087 -663
rect 2029 -731 2087 -697
rect 2029 -765 2041 -731
rect 2075 -765 2087 -731
rect 2029 -799 2087 -765
rect 2029 -833 2041 -799
rect 2075 -833 2087 -799
rect 2029 -867 2087 -833
rect 2029 -901 2041 -867
rect 2075 -901 2087 -867
rect 2029 -935 2087 -901
rect 2029 -969 2041 -935
rect 2075 -969 2087 -935
rect 2029 -1003 2087 -969
rect 2029 -1037 2041 -1003
rect 2075 -1037 2087 -1003
rect 2029 -1071 2087 -1037
rect 2029 -1105 2041 -1071
rect 2075 -1105 2087 -1071
rect 2029 -1139 2087 -1105
rect 2029 -1173 2041 -1139
rect 2075 -1173 2087 -1139
rect 2029 -1207 2087 -1173
rect 2029 -1241 2041 -1207
rect 2075 -1241 2087 -1207
rect 2029 -1275 2087 -1241
rect 2029 -1309 2041 -1275
rect 2075 -1309 2087 -1275
rect 2029 -1343 2087 -1309
rect 2029 -1377 2041 -1343
rect 2075 -1377 2087 -1343
rect 2029 -1411 2087 -1377
rect 2029 -1445 2041 -1411
rect 2075 -1445 2087 -1411
rect 2029 -1479 2087 -1445
rect 2029 -1513 2041 -1479
rect 2075 -1513 2087 -1479
rect 2029 -1547 2087 -1513
rect 2029 -1581 2041 -1547
rect 2075 -1581 2087 -1547
rect 2029 -1615 2087 -1581
rect 2029 -1649 2041 -1615
rect 2075 -1649 2087 -1615
rect 2029 -1683 2087 -1649
rect 2029 -1717 2041 -1683
rect 2075 -1717 2087 -1683
rect 2029 -1751 2087 -1717
rect 2029 -1785 2041 -1751
rect 2075 -1785 2087 -1751
rect 2029 -1819 2087 -1785
rect 2029 -1853 2041 -1819
rect 2075 -1853 2087 -1819
rect 2029 -1887 2087 -1853
rect 2029 -1921 2041 -1887
rect 2075 -1921 2087 -1887
rect 2029 -1955 2087 -1921
rect 2029 -1989 2041 -1955
rect 2075 -1989 2087 -1955
rect 2029 -2023 2087 -1989
rect 2029 -2057 2041 -2023
rect 2075 -2057 2087 -2023
rect 2029 -2091 2087 -2057
rect 2029 -2125 2041 -2091
rect 2075 -2125 2087 -2091
rect 2029 -2159 2087 -2125
rect 2029 -2193 2041 -2159
rect 2075 -2193 2087 -2159
rect 2029 -2227 2087 -2193
rect 2029 -2261 2041 -2227
rect 2075 -2261 2087 -2227
rect 2029 -2295 2087 -2261
rect 2029 -2329 2041 -2295
rect 2075 -2329 2087 -2295
rect 2029 -2363 2087 -2329
rect 2029 -2397 2041 -2363
rect 2075 -2397 2087 -2363
rect 2029 -2431 2087 -2397
rect 2029 -2465 2041 -2431
rect 2075 -2465 2087 -2431
rect 2029 -2500 2087 -2465
rect 4087 2465 4145 2500
rect 4087 2431 4099 2465
rect 4133 2431 4145 2465
rect 4087 2397 4145 2431
rect 4087 2363 4099 2397
rect 4133 2363 4145 2397
rect 4087 2329 4145 2363
rect 4087 2295 4099 2329
rect 4133 2295 4145 2329
rect 4087 2261 4145 2295
rect 4087 2227 4099 2261
rect 4133 2227 4145 2261
rect 4087 2193 4145 2227
rect 4087 2159 4099 2193
rect 4133 2159 4145 2193
rect 4087 2125 4145 2159
rect 4087 2091 4099 2125
rect 4133 2091 4145 2125
rect 4087 2057 4145 2091
rect 4087 2023 4099 2057
rect 4133 2023 4145 2057
rect 4087 1989 4145 2023
rect 4087 1955 4099 1989
rect 4133 1955 4145 1989
rect 4087 1921 4145 1955
rect 4087 1887 4099 1921
rect 4133 1887 4145 1921
rect 4087 1853 4145 1887
rect 4087 1819 4099 1853
rect 4133 1819 4145 1853
rect 4087 1785 4145 1819
rect 4087 1751 4099 1785
rect 4133 1751 4145 1785
rect 4087 1717 4145 1751
rect 4087 1683 4099 1717
rect 4133 1683 4145 1717
rect 4087 1649 4145 1683
rect 4087 1615 4099 1649
rect 4133 1615 4145 1649
rect 4087 1581 4145 1615
rect 4087 1547 4099 1581
rect 4133 1547 4145 1581
rect 4087 1513 4145 1547
rect 4087 1479 4099 1513
rect 4133 1479 4145 1513
rect 4087 1445 4145 1479
rect 4087 1411 4099 1445
rect 4133 1411 4145 1445
rect 4087 1377 4145 1411
rect 4087 1343 4099 1377
rect 4133 1343 4145 1377
rect 4087 1309 4145 1343
rect 4087 1275 4099 1309
rect 4133 1275 4145 1309
rect 4087 1241 4145 1275
rect 4087 1207 4099 1241
rect 4133 1207 4145 1241
rect 4087 1173 4145 1207
rect 4087 1139 4099 1173
rect 4133 1139 4145 1173
rect 4087 1105 4145 1139
rect 4087 1071 4099 1105
rect 4133 1071 4145 1105
rect 4087 1037 4145 1071
rect 4087 1003 4099 1037
rect 4133 1003 4145 1037
rect 4087 969 4145 1003
rect 4087 935 4099 969
rect 4133 935 4145 969
rect 4087 901 4145 935
rect 4087 867 4099 901
rect 4133 867 4145 901
rect 4087 833 4145 867
rect 4087 799 4099 833
rect 4133 799 4145 833
rect 4087 765 4145 799
rect 4087 731 4099 765
rect 4133 731 4145 765
rect 4087 697 4145 731
rect 4087 663 4099 697
rect 4133 663 4145 697
rect 4087 629 4145 663
rect 4087 595 4099 629
rect 4133 595 4145 629
rect 4087 561 4145 595
rect 4087 527 4099 561
rect 4133 527 4145 561
rect 4087 493 4145 527
rect 4087 459 4099 493
rect 4133 459 4145 493
rect 4087 425 4145 459
rect 4087 391 4099 425
rect 4133 391 4145 425
rect 4087 357 4145 391
rect 4087 323 4099 357
rect 4133 323 4145 357
rect 4087 289 4145 323
rect 4087 255 4099 289
rect 4133 255 4145 289
rect 4087 221 4145 255
rect 4087 187 4099 221
rect 4133 187 4145 221
rect 4087 153 4145 187
rect 4087 119 4099 153
rect 4133 119 4145 153
rect 4087 85 4145 119
rect 4087 51 4099 85
rect 4133 51 4145 85
rect 4087 17 4145 51
rect 4087 -17 4099 17
rect 4133 -17 4145 17
rect 4087 -51 4145 -17
rect 4087 -85 4099 -51
rect 4133 -85 4145 -51
rect 4087 -119 4145 -85
rect 4087 -153 4099 -119
rect 4133 -153 4145 -119
rect 4087 -187 4145 -153
rect 4087 -221 4099 -187
rect 4133 -221 4145 -187
rect 4087 -255 4145 -221
rect 4087 -289 4099 -255
rect 4133 -289 4145 -255
rect 4087 -323 4145 -289
rect 4087 -357 4099 -323
rect 4133 -357 4145 -323
rect 4087 -391 4145 -357
rect 4087 -425 4099 -391
rect 4133 -425 4145 -391
rect 4087 -459 4145 -425
rect 4087 -493 4099 -459
rect 4133 -493 4145 -459
rect 4087 -527 4145 -493
rect 4087 -561 4099 -527
rect 4133 -561 4145 -527
rect 4087 -595 4145 -561
rect 4087 -629 4099 -595
rect 4133 -629 4145 -595
rect 4087 -663 4145 -629
rect 4087 -697 4099 -663
rect 4133 -697 4145 -663
rect 4087 -731 4145 -697
rect 4087 -765 4099 -731
rect 4133 -765 4145 -731
rect 4087 -799 4145 -765
rect 4087 -833 4099 -799
rect 4133 -833 4145 -799
rect 4087 -867 4145 -833
rect 4087 -901 4099 -867
rect 4133 -901 4145 -867
rect 4087 -935 4145 -901
rect 4087 -969 4099 -935
rect 4133 -969 4145 -935
rect 4087 -1003 4145 -969
rect 4087 -1037 4099 -1003
rect 4133 -1037 4145 -1003
rect 4087 -1071 4145 -1037
rect 4087 -1105 4099 -1071
rect 4133 -1105 4145 -1071
rect 4087 -1139 4145 -1105
rect 4087 -1173 4099 -1139
rect 4133 -1173 4145 -1139
rect 4087 -1207 4145 -1173
rect 4087 -1241 4099 -1207
rect 4133 -1241 4145 -1207
rect 4087 -1275 4145 -1241
rect 4087 -1309 4099 -1275
rect 4133 -1309 4145 -1275
rect 4087 -1343 4145 -1309
rect 4087 -1377 4099 -1343
rect 4133 -1377 4145 -1343
rect 4087 -1411 4145 -1377
rect 4087 -1445 4099 -1411
rect 4133 -1445 4145 -1411
rect 4087 -1479 4145 -1445
rect 4087 -1513 4099 -1479
rect 4133 -1513 4145 -1479
rect 4087 -1547 4145 -1513
rect 4087 -1581 4099 -1547
rect 4133 -1581 4145 -1547
rect 4087 -1615 4145 -1581
rect 4087 -1649 4099 -1615
rect 4133 -1649 4145 -1615
rect 4087 -1683 4145 -1649
rect 4087 -1717 4099 -1683
rect 4133 -1717 4145 -1683
rect 4087 -1751 4145 -1717
rect 4087 -1785 4099 -1751
rect 4133 -1785 4145 -1751
rect 4087 -1819 4145 -1785
rect 4087 -1853 4099 -1819
rect 4133 -1853 4145 -1819
rect 4087 -1887 4145 -1853
rect 4087 -1921 4099 -1887
rect 4133 -1921 4145 -1887
rect 4087 -1955 4145 -1921
rect 4087 -1989 4099 -1955
rect 4133 -1989 4145 -1955
rect 4087 -2023 4145 -1989
rect 4087 -2057 4099 -2023
rect 4133 -2057 4145 -2023
rect 4087 -2091 4145 -2057
rect 4087 -2125 4099 -2091
rect 4133 -2125 4145 -2091
rect 4087 -2159 4145 -2125
rect 4087 -2193 4099 -2159
rect 4133 -2193 4145 -2159
rect 4087 -2227 4145 -2193
rect 4087 -2261 4099 -2227
rect 4133 -2261 4145 -2227
rect 4087 -2295 4145 -2261
rect 4087 -2329 4099 -2295
rect 4133 -2329 4145 -2295
rect 4087 -2363 4145 -2329
rect 4087 -2397 4099 -2363
rect 4133 -2397 4145 -2363
rect 4087 -2431 4145 -2397
rect 4087 -2465 4099 -2431
rect 4133 -2465 4145 -2431
rect 4087 -2500 4145 -2465
<< ndiffc >>
rect -4133 2431 -4099 2465
rect -4133 2363 -4099 2397
rect -4133 2295 -4099 2329
rect -4133 2227 -4099 2261
rect -4133 2159 -4099 2193
rect -4133 2091 -4099 2125
rect -4133 2023 -4099 2057
rect -4133 1955 -4099 1989
rect -4133 1887 -4099 1921
rect -4133 1819 -4099 1853
rect -4133 1751 -4099 1785
rect -4133 1683 -4099 1717
rect -4133 1615 -4099 1649
rect -4133 1547 -4099 1581
rect -4133 1479 -4099 1513
rect -4133 1411 -4099 1445
rect -4133 1343 -4099 1377
rect -4133 1275 -4099 1309
rect -4133 1207 -4099 1241
rect -4133 1139 -4099 1173
rect -4133 1071 -4099 1105
rect -4133 1003 -4099 1037
rect -4133 935 -4099 969
rect -4133 867 -4099 901
rect -4133 799 -4099 833
rect -4133 731 -4099 765
rect -4133 663 -4099 697
rect -4133 595 -4099 629
rect -4133 527 -4099 561
rect -4133 459 -4099 493
rect -4133 391 -4099 425
rect -4133 323 -4099 357
rect -4133 255 -4099 289
rect -4133 187 -4099 221
rect -4133 119 -4099 153
rect -4133 51 -4099 85
rect -4133 -17 -4099 17
rect -4133 -85 -4099 -51
rect -4133 -153 -4099 -119
rect -4133 -221 -4099 -187
rect -4133 -289 -4099 -255
rect -4133 -357 -4099 -323
rect -4133 -425 -4099 -391
rect -4133 -493 -4099 -459
rect -4133 -561 -4099 -527
rect -4133 -629 -4099 -595
rect -4133 -697 -4099 -663
rect -4133 -765 -4099 -731
rect -4133 -833 -4099 -799
rect -4133 -901 -4099 -867
rect -4133 -969 -4099 -935
rect -4133 -1037 -4099 -1003
rect -4133 -1105 -4099 -1071
rect -4133 -1173 -4099 -1139
rect -4133 -1241 -4099 -1207
rect -4133 -1309 -4099 -1275
rect -4133 -1377 -4099 -1343
rect -4133 -1445 -4099 -1411
rect -4133 -1513 -4099 -1479
rect -4133 -1581 -4099 -1547
rect -4133 -1649 -4099 -1615
rect -4133 -1717 -4099 -1683
rect -4133 -1785 -4099 -1751
rect -4133 -1853 -4099 -1819
rect -4133 -1921 -4099 -1887
rect -4133 -1989 -4099 -1955
rect -4133 -2057 -4099 -2023
rect -4133 -2125 -4099 -2091
rect -4133 -2193 -4099 -2159
rect -4133 -2261 -4099 -2227
rect -4133 -2329 -4099 -2295
rect -4133 -2397 -4099 -2363
rect -4133 -2465 -4099 -2431
rect -2075 2431 -2041 2465
rect -2075 2363 -2041 2397
rect -2075 2295 -2041 2329
rect -2075 2227 -2041 2261
rect -2075 2159 -2041 2193
rect -2075 2091 -2041 2125
rect -2075 2023 -2041 2057
rect -2075 1955 -2041 1989
rect -2075 1887 -2041 1921
rect -2075 1819 -2041 1853
rect -2075 1751 -2041 1785
rect -2075 1683 -2041 1717
rect -2075 1615 -2041 1649
rect -2075 1547 -2041 1581
rect -2075 1479 -2041 1513
rect -2075 1411 -2041 1445
rect -2075 1343 -2041 1377
rect -2075 1275 -2041 1309
rect -2075 1207 -2041 1241
rect -2075 1139 -2041 1173
rect -2075 1071 -2041 1105
rect -2075 1003 -2041 1037
rect -2075 935 -2041 969
rect -2075 867 -2041 901
rect -2075 799 -2041 833
rect -2075 731 -2041 765
rect -2075 663 -2041 697
rect -2075 595 -2041 629
rect -2075 527 -2041 561
rect -2075 459 -2041 493
rect -2075 391 -2041 425
rect -2075 323 -2041 357
rect -2075 255 -2041 289
rect -2075 187 -2041 221
rect -2075 119 -2041 153
rect -2075 51 -2041 85
rect -2075 -17 -2041 17
rect -2075 -85 -2041 -51
rect -2075 -153 -2041 -119
rect -2075 -221 -2041 -187
rect -2075 -289 -2041 -255
rect -2075 -357 -2041 -323
rect -2075 -425 -2041 -391
rect -2075 -493 -2041 -459
rect -2075 -561 -2041 -527
rect -2075 -629 -2041 -595
rect -2075 -697 -2041 -663
rect -2075 -765 -2041 -731
rect -2075 -833 -2041 -799
rect -2075 -901 -2041 -867
rect -2075 -969 -2041 -935
rect -2075 -1037 -2041 -1003
rect -2075 -1105 -2041 -1071
rect -2075 -1173 -2041 -1139
rect -2075 -1241 -2041 -1207
rect -2075 -1309 -2041 -1275
rect -2075 -1377 -2041 -1343
rect -2075 -1445 -2041 -1411
rect -2075 -1513 -2041 -1479
rect -2075 -1581 -2041 -1547
rect -2075 -1649 -2041 -1615
rect -2075 -1717 -2041 -1683
rect -2075 -1785 -2041 -1751
rect -2075 -1853 -2041 -1819
rect -2075 -1921 -2041 -1887
rect -2075 -1989 -2041 -1955
rect -2075 -2057 -2041 -2023
rect -2075 -2125 -2041 -2091
rect -2075 -2193 -2041 -2159
rect -2075 -2261 -2041 -2227
rect -2075 -2329 -2041 -2295
rect -2075 -2397 -2041 -2363
rect -2075 -2465 -2041 -2431
rect -17 2431 17 2465
rect -17 2363 17 2397
rect -17 2295 17 2329
rect -17 2227 17 2261
rect -17 2159 17 2193
rect -17 2091 17 2125
rect -17 2023 17 2057
rect -17 1955 17 1989
rect -17 1887 17 1921
rect -17 1819 17 1853
rect -17 1751 17 1785
rect -17 1683 17 1717
rect -17 1615 17 1649
rect -17 1547 17 1581
rect -17 1479 17 1513
rect -17 1411 17 1445
rect -17 1343 17 1377
rect -17 1275 17 1309
rect -17 1207 17 1241
rect -17 1139 17 1173
rect -17 1071 17 1105
rect -17 1003 17 1037
rect -17 935 17 969
rect -17 867 17 901
rect -17 799 17 833
rect -17 731 17 765
rect -17 663 17 697
rect -17 595 17 629
rect -17 527 17 561
rect -17 459 17 493
rect -17 391 17 425
rect -17 323 17 357
rect -17 255 17 289
rect -17 187 17 221
rect -17 119 17 153
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect -17 -153 17 -119
rect -17 -221 17 -187
rect -17 -289 17 -255
rect -17 -357 17 -323
rect -17 -425 17 -391
rect -17 -493 17 -459
rect -17 -561 17 -527
rect -17 -629 17 -595
rect -17 -697 17 -663
rect -17 -765 17 -731
rect -17 -833 17 -799
rect -17 -901 17 -867
rect -17 -969 17 -935
rect -17 -1037 17 -1003
rect -17 -1105 17 -1071
rect -17 -1173 17 -1139
rect -17 -1241 17 -1207
rect -17 -1309 17 -1275
rect -17 -1377 17 -1343
rect -17 -1445 17 -1411
rect -17 -1513 17 -1479
rect -17 -1581 17 -1547
rect -17 -1649 17 -1615
rect -17 -1717 17 -1683
rect -17 -1785 17 -1751
rect -17 -1853 17 -1819
rect -17 -1921 17 -1887
rect -17 -1989 17 -1955
rect -17 -2057 17 -2023
rect -17 -2125 17 -2091
rect -17 -2193 17 -2159
rect -17 -2261 17 -2227
rect -17 -2329 17 -2295
rect -17 -2397 17 -2363
rect -17 -2465 17 -2431
rect 2041 2431 2075 2465
rect 2041 2363 2075 2397
rect 2041 2295 2075 2329
rect 2041 2227 2075 2261
rect 2041 2159 2075 2193
rect 2041 2091 2075 2125
rect 2041 2023 2075 2057
rect 2041 1955 2075 1989
rect 2041 1887 2075 1921
rect 2041 1819 2075 1853
rect 2041 1751 2075 1785
rect 2041 1683 2075 1717
rect 2041 1615 2075 1649
rect 2041 1547 2075 1581
rect 2041 1479 2075 1513
rect 2041 1411 2075 1445
rect 2041 1343 2075 1377
rect 2041 1275 2075 1309
rect 2041 1207 2075 1241
rect 2041 1139 2075 1173
rect 2041 1071 2075 1105
rect 2041 1003 2075 1037
rect 2041 935 2075 969
rect 2041 867 2075 901
rect 2041 799 2075 833
rect 2041 731 2075 765
rect 2041 663 2075 697
rect 2041 595 2075 629
rect 2041 527 2075 561
rect 2041 459 2075 493
rect 2041 391 2075 425
rect 2041 323 2075 357
rect 2041 255 2075 289
rect 2041 187 2075 221
rect 2041 119 2075 153
rect 2041 51 2075 85
rect 2041 -17 2075 17
rect 2041 -85 2075 -51
rect 2041 -153 2075 -119
rect 2041 -221 2075 -187
rect 2041 -289 2075 -255
rect 2041 -357 2075 -323
rect 2041 -425 2075 -391
rect 2041 -493 2075 -459
rect 2041 -561 2075 -527
rect 2041 -629 2075 -595
rect 2041 -697 2075 -663
rect 2041 -765 2075 -731
rect 2041 -833 2075 -799
rect 2041 -901 2075 -867
rect 2041 -969 2075 -935
rect 2041 -1037 2075 -1003
rect 2041 -1105 2075 -1071
rect 2041 -1173 2075 -1139
rect 2041 -1241 2075 -1207
rect 2041 -1309 2075 -1275
rect 2041 -1377 2075 -1343
rect 2041 -1445 2075 -1411
rect 2041 -1513 2075 -1479
rect 2041 -1581 2075 -1547
rect 2041 -1649 2075 -1615
rect 2041 -1717 2075 -1683
rect 2041 -1785 2075 -1751
rect 2041 -1853 2075 -1819
rect 2041 -1921 2075 -1887
rect 2041 -1989 2075 -1955
rect 2041 -2057 2075 -2023
rect 2041 -2125 2075 -2091
rect 2041 -2193 2075 -2159
rect 2041 -2261 2075 -2227
rect 2041 -2329 2075 -2295
rect 2041 -2397 2075 -2363
rect 2041 -2465 2075 -2431
rect 4099 2431 4133 2465
rect 4099 2363 4133 2397
rect 4099 2295 4133 2329
rect 4099 2227 4133 2261
rect 4099 2159 4133 2193
rect 4099 2091 4133 2125
rect 4099 2023 4133 2057
rect 4099 1955 4133 1989
rect 4099 1887 4133 1921
rect 4099 1819 4133 1853
rect 4099 1751 4133 1785
rect 4099 1683 4133 1717
rect 4099 1615 4133 1649
rect 4099 1547 4133 1581
rect 4099 1479 4133 1513
rect 4099 1411 4133 1445
rect 4099 1343 4133 1377
rect 4099 1275 4133 1309
rect 4099 1207 4133 1241
rect 4099 1139 4133 1173
rect 4099 1071 4133 1105
rect 4099 1003 4133 1037
rect 4099 935 4133 969
rect 4099 867 4133 901
rect 4099 799 4133 833
rect 4099 731 4133 765
rect 4099 663 4133 697
rect 4099 595 4133 629
rect 4099 527 4133 561
rect 4099 459 4133 493
rect 4099 391 4133 425
rect 4099 323 4133 357
rect 4099 255 4133 289
rect 4099 187 4133 221
rect 4099 119 4133 153
rect 4099 51 4133 85
rect 4099 -17 4133 17
rect 4099 -85 4133 -51
rect 4099 -153 4133 -119
rect 4099 -221 4133 -187
rect 4099 -289 4133 -255
rect 4099 -357 4133 -323
rect 4099 -425 4133 -391
rect 4099 -493 4133 -459
rect 4099 -561 4133 -527
rect 4099 -629 4133 -595
rect 4099 -697 4133 -663
rect 4099 -765 4133 -731
rect 4099 -833 4133 -799
rect 4099 -901 4133 -867
rect 4099 -969 4133 -935
rect 4099 -1037 4133 -1003
rect 4099 -1105 4133 -1071
rect 4099 -1173 4133 -1139
rect 4099 -1241 4133 -1207
rect 4099 -1309 4133 -1275
rect 4099 -1377 4133 -1343
rect 4099 -1445 4133 -1411
rect 4099 -1513 4133 -1479
rect 4099 -1581 4133 -1547
rect 4099 -1649 4133 -1615
rect 4099 -1717 4133 -1683
rect 4099 -1785 4133 -1751
rect 4099 -1853 4133 -1819
rect 4099 -1921 4133 -1887
rect 4099 -1989 4133 -1955
rect 4099 -2057 4133 -2023
rect 4099 -2125 4133 -2091
rect 4099 -2193 4133 -2159
rect 4099 -2261 4133 -2227
rect 4099 -2329 4133 -2295
rect 4099 -2397 4133 -2363
rect 4099 -2465 4133 -2431
<< psubdiff >>
rect -4247 2640 -4131 2674
rect -4097 2640 -4063 2674
rect -4029 2640 -3995 2674
rect -3961 2640 -3927 2674
rect -3893 2640 -3859 2674
rect -3825 2640 -3791 2674
rect -3757 2640 -3723 2674
rect -3689 2640 -3655 2674
rect -3621 2640 -3587 2674
rect -3553 2640 -3519 2674
rect -3485 2640 -3451 2674
rect -3417 2640 -3383 2674
rect -3349 2640 -3315 2674
rect -3281 2640 -3247 2674
rect -3213 2640 -3179 2674
rect -3145 2640 -3111 2674
rect -3077 2640 -3043 2674
rect -3009 2640 -2975 2674
rect -2941 2640 -2907 2674
rect -2873 2640 -2839 2674
rect -2805 2640 -2771 2674
rect -2737 2640 -2703 2674
rect -2669 2640 -2635 2674
rect -2601 2640 -2567 2674
rect -2533 2640 -2499 2674
rect -2465 2640 -2431 2674
rect -2397 2640 -2363 2674
rect -2329 2640 -2295 2674
rect -2261 2640 -2227 2674
rect -2193 2640 -2159 2674
rect -2125 2640 -2091 2674
rect -2057 2640 -2023 2674
rect -1989 2640 -1955 2674
rect -1921 2640 -1887 2674
rect -1853 2640 -1819 2674
rect -1785 2640 -1751 2674
rect -1717 2640 -1683 2674
rect -1649 2640 -1615 2674
rect -1581 2640 -1547 2674
rect -1513 2640 -1479 2674
rect -1445 2640 -1411 2674
rect -1377 2640 -1343 2674
rect -1309 2640 -1275 2674
rect -1241 2640 -1207 2674
rect -1173 2640 -1139 2674
rect -1105 2640 -1071 2674
rect -1037 2640 -1003 2674
rect -969 2640 -935 2674
rect -901 2640 -867 2674
rect -833 2640 -799 2674
rect -765 2640 -731 2674
rect -697 2640 -663 2674
rect -629 2640 -595 2674
rect -561 2640 -527 2674
rect -493 2640 -459 2674
rect -425 2640 -391 2674
rect -357 2640 -323 2674
rect -289 2640 -255 2674
rect -221 2640 -187 2674
rect -153 2640 -119 2674
rect -85 2640 -51 2674
rect -17 2640 17 2674
rect 51 2640 85 2674
rect 119 2640 153 2674
rect 187 2640 221 2674
rect 255 2640 289 2674
rect 323 2640 357 2674
rect 391 2640 425 2674
rect 459 2640 493 2674
rect 527 2640 561 2674
rect 595 2640 629 2674
rect 663 2640 697 2674
rect 731 2640 765 2674
rect 799 2640 833 2674
rect 867 2640 901 2674
rect 935 2640 969 2674
rect 1003 2640 1037 2674
rect 1071 2640 1105 2674
rect 1139 2640 1173 2674
rect 1207 2640 1241 2674
rect 1275 2640 1309 2674
rect 1343 2640 1377 2674
rect 1411 2640 1445 2674
rect 1479 2640 1513 2674
rect 1547 2640 1581 2674
rect 1615 2640 1649 2674
rect 1683 2640 1717 2674
rect 1751 2640 1785 2674
rect 1819 2640 1853 2674
rect 1887 2640 1921 2674
rect 1955 2640 1989 2674
rect 2023 2640 2057 2674
rect 2091 2640 2125 2674
rect 2159 2640 2193 2674
rect 2227 2640 2261 2674
rect 2295 2640 2329 2674
rect 2363 2640 2397 2674
rect 2431 2640 2465 2674
rect 2499 2640 2533 2674
rect 2567 2640 2601 2674
rect 2635 2640 2669 2674
rect 2703 2640 2737 2674
rect 2771 2640 2805 2674
rect 2839 2640 2873 2674
rect 2907 2640 2941 2674
rect 2975 2640 3009 2674
rect 3043 2640 3077 2674
rect 3111 2640 3145 2674
rect 3179 2640 3213 2674
rect 3247 2640 3281 2674
rect 3315 2640 3349 2674
rect 3383 2640 3417 2674
rect 3451 2640 3485 2674
rect 3519 2640 3553 2674
rect 3587 2640 3621 2674
rect 3655 2640 3689 2674
rect 3723 2640 3757 2674
rect 3791 2640 3825 2674
rect 3859 2640 3893 2674
rect 3927 2640 3961 2674
rect 3995 2640 4029 2674
rect 4063 2640 4097 2674
rect 4131 2640 4247 2674
rect -4247 2567 -4213 2640
rect -4247 2499 -4213 2533
rect 4213 2567 4247 2640
rect -4247 2431 -4213 2465
rect -4247 2363 -4213 2397
rect -4247 2295 -4213 2329
rect -4247 2227 -4213 2261
rect -4247 2159 -4213 2193
rect -4247 2091 -4213 2125
rect -4247 2023 -4213 2057
rect -4247 1955 -4213 1989
rect -4247 1887 -4213 1921
rect -4247 1819 -4213 1853
rect -4247 1751 -4213 1785
rect -4247 1683 -4213 1717
rect -4247 1615 -4213 1649
rect -4247 1547 -4213 1581
rect -4247 1479 -4213 1513
rect -4247 1411 -4213 1445
rect -4247 1343 -4213 1377
rect -4247 1275 -4213 1309
rect -4247 1207 -4213 1241
rect -4247 1139 -4213 1173
rect -4247 1071 -4213 1105
rect -4247 1003 -4213 1037
rect -4247 935 -4213 969
rect -4247 867 -4213 901
rect -4247 799 -4213 833
rect -4247 731 -4213 765
rect -4247 663 -4213 697
rect -4247 595 -4213 629
rect -4247 527 -4213 561
rect -4247 459 -4213 493
rect -4247 391 -4213 425
rect -4247 323 -4213 357
rect -4247 255 -4213 289
rect -4247 187 -4213 221
rect -4247 119 -4213 153
rect -4247 51 -4213 85
rect -4247 -17 -4213 17
rect -4247 -85 -4213 -51
rect -4247 -153 -4213 -119
rect -4247 -221 -4213 -187
rect -4247 -289 -4213 -255
rect -4247 -357 -4213 -323
rect -4247 -425 -4213 -391
rect -4247 -493 -4213 -459
rect -4247 -561 -4213 -527
rect -4247 -629 -4213 -595
rect -4247 -697 -4213 -663
rect -4247 -765 -4213 -731
rect -4247 -833 -4213 -799
rect -4247 -901 -4213 -867
rect -4247 -969 -4213 -935
rect -4247 -1037 -4213 -1003
rect -4247 -1105 -4213 -1071
rect -4247 -1173 -4213 -1139
rect -4247 -1241 -4213 -1207
rect -4247 -1309 -4213 -1275
rect -4247 -1377 -4213 -1343
rect -4247 -1445 -4213 -1411
rect -4247 -1513 -4213 -1479
rect -4247 -1581 -4213 -1547
rect -4247 -1649 -4213 -1615
rect -4247 -1717 -4213 -1683
rect -4247 -1785 -4213 -1751
rect -4247 -1853 -4213 -1819
rect -4247 -1921 -4213 -1887
rect -4247 -1989 -4213 -1955
rect -4247 -2057 -4213 -2023
rect -4247 -2125 -4213 -2091
rect -4247 -2193 -4213 -2159
rect -4247 -2261 -4213 -2227
rect -4247 -2329 -4213 -2295
rect -4247 -2397 -4213 -2363
rect -4247 -2465 -4213 -2431
rect -4247 -2533 -4213 -2499
rect 4213 2499 4247 2533
rect 4213 2431 4247 2465
rect 4213 2363 4247 2397
rect 4213 2295 4247 2329
rect 4213 2227 4247 2261
rect 4213 2159 4247 2193
rect 4213 2091 4247 2125
rect 4213 2023 4247 2057
rect 4213 1955 4247 1989
rect 4213 1887 4247 1921
rect 4213 1819 4247 1853
rect 4213 1751 4247 1785
rect 4213 1683 4247 1717
rect 4213 1615 4247 1649
rect 4213 1547 4247 1581
rect 4213 1479 4247 1513
rect 4213 1411 4247 1445
rect 4213 1343 4247 1377
rect 4213 1275 4247 1309
rect 4213 1207 4247 1241
rect 4213 1139 4247 1173
rect 4213 1071 4247 1105
rect 4213 1003 4247 1037
rect 4213 935 4247 969
rect 4213 867 4247 901
rect 4213 799 4247 833
rect 4213 731 4247 765
rect 4213 663 4247 697
rect 4213 595 4247 629
rect 4213 527 4247 561
rect 4213 459 4247 493
rect 4213 391 4247 425
rect 4213 323 4247 357
rect 4213 255 4247 289
rect 4213 187 4247 221
rect 4213 119 4247 153
rect 4213 51 4247 85
rect 4213 -17 4247 17
rect 4213 -85 4247 -51
rect 4213 -153 4247 -119
rect 4213 -221 4247 -187
rect 4213 -289 4247 -255
rect 4213 -357 4247 -323
rect 4213 -425 4247 -391
rect 4213 -493 4247 -459
rect 4213 -561 4247 -527
rect 4213 -629 4247 -595
rect 4213 -697 4247 -663
rect 4213 -765 4247 -731
rect 4213 -833 4247 -799
rect 4213 -901 4247 -867
rect 4213 -969 4247 -935
rect 4213 -1037 4247 -1003
rect 4213 -1105 4247 -1071
rect 4213 -1173 4247 -1139
rect 4213 -1241 4247 -1207
rect 4213 -1309 4247 -1275
rect 4213 -1377 4247 -1343
rect 4213 -1445 4247 -1411
rect 4213 -1513 4247 -1479
rect 4213 -1581 4247 -1547
rect 4213 -1649 4247 -1615
rect 4213 -1717 4247 -1683
rect 4213 -1785 4247 -1751
rect 4213 -1853 4247 -1819
rect 4213 -1921 4247 -1887
rect 4213 -1989 4247 -1955
rect 4213 -2057 4247 -2023
rect 4213 -2125 4247 -2091
rect 4213 -2193 4247 -2159
rect 4213 -2261 4247 -2227
rect 4213 -2329 4247 -2295
rect 4213 -2397 4247 -2363
rect 4213 -2465 4247 -2431
rect -4247 -2640 -4213 -2567
rect 4213 -2533 4247 -2499
rect 4213 -2640 4247 -2567
rect -4247 -2674 -4131 -2640
rect -4097 -2674 -4063 -2640
rect -4029 -2674 -3995 -2640
rect -3961 -2674 -3927 -2640
rect -3893 -2674 -3859 -2640
rect -3825 -2674 -3791 -2640
rect -3757 -2674 -3723 -2640
rect -3689 -2674 -3655 -2640
rect -3621 -2674 -3587 -2640
rect -3553 -2674 -3519 -2640
rect -3485 -2674 -3451 -2640
rect -3417 -2674 -3383 -2640
rect -3349 -2674 -3315 -2640
rect -3281 -2674 -3247 -2640
rect -3213 -2674 -3179 -2640
rect -3145 -2674 -3111 -2640
rect -3077 -2674 -3043 -2640
rect -3009 -2674 -2975 -2640
rect -2941 -2674 -2907 -2640
rect -2873 -2674 -2839 -2640
rect -2805 -2674 -2771 -2640
rect -2737 -2674 -2703 -2640
rect -2669 -2674 -2635 -2640
rect -2601 -2674 -2567 -2640
rect -2533 -2674 -2499 -2640
rect -2465 -2674 -2431 -2640
rect -2397 -2674 -2363 -2640
rect -2329 -2674 -2295 -2640
rect -2261 -2674 -2227 -2640
rect -2193 -2674 -2159 -2640
rect -2125 -2674 -2091 -2640
rect -2057 -2674 -2023 -2640
rect -1989 -2674 -1955 -2640
rect -1921 -2674 -1887 -2640
rect -1853 -2674 -1819 -2640
rect -1785 -2674 -1751 -2640
rect -1717 -2674 -1683 -2640
rect -1649 -2674 -1615 -2640
rect -1581 -2674 -1547 -2640
rect -1513 -2674 -1479 -2640
rect -1445 -2674 -1411 -2640
rect -1377 -2674 -1343 -2640
rect -1309 -2674 -1275 -2640
rect -1241 -2674 -1207 -2640
rect -1173 -2674 -1139 -2640
rect -1105 -2674 -1071 -2640
rect -1037 -2674 -1003 -2640
rect -969 -2674 -935 -2640
rect -901 -2674 -867 -2640
rect -833 -2674 -799 -2640
rect -765 -2674 -731 -2640
rect -697 -2674 -663 -2640
rect -629 -2674 -595 -2640
rect -561 -2674 -527 -2640
rect -493 -2674 -459 -2640
rect -425 -2674 -391 -2640
rect -357 -2674 -323 -2640
rect -289 -2674 -255 -2640
rect -221 -2674 -187 -2640
rect -153 -2674 -119 -2640
rect -85 -2674 -51 -2640
rect -17 -2674 17 -2640
rect 51 -2674 85 -2640
rect 119 -2674 153 -2640
rect 187 -2674 221 -2640
rect 255 -2674 289 -2640
rect 323 -2674 357 -2640
rect 391 -2674 425 -2640
rect 459 -2674 493 -2640
rect 527 -2674 561 -2640
rect 595 -2674 629 -2640
rect 663 -2674 697 -2640
rect 731 -2674 765 -2640
rect 799 -2674 833 -2640
rect 867 -2674 901 -2640
rect 935 -2674 969 -2640
rect 1003 -2674 1037 -2640
rect 1071 -2674 1105 -2640
rect 1139 -2674 1173 -2640
rect 1207 -2674 1241 -2640
rect 1275 -2674 1309 -2640
rect 1343 -2674 1377 -2640
rect 1411 -2674 1445 -2640
rect 1479 -2674 1513 -2640
rect 1547 -2674 1581 -2640
rect 1615 -2674 1649 -2640
rect 1683 -2674 1717 -2640
rect 1751 -2674 1785 -2640
rect 1819 -2674 1853 -2640
rect 1887 -2674 1921 -2640
rect 1955 -2674 1989 -2640
rect 2023 -2674 2057 -2640
rect 2091 -2674 2125 -2640
rect 2159 -2674 2193 -2640
rect 2227 -2674 2261 -2640
rect 2295 -2674 2329 -2640
rect 2363 -2674 2397 -2640
rect 2431 -2674 2465 -2640
rect 2499 -2674 2533 -2640
rect 2567 -2674 2601 -2640
rect 2635 -2674 2669 -2640
rect 2703 -2674 2737 -2640
rect 2771 -2674 2805 -2640
rect 2839 -2674 2873 -2640
rect 2907 -2674 2941 -2640
rect 2975 -2674 3009 -2640
rect 3043 -2674 3077 -2640
rect 3111 -2674 3145 -2640
rect 3179 -2674 3213 -2640
rect 3247 -2674 3281 -2640
rect 3315 -2674 3349 -2640
rect 3383 -2674 3417 -2640
rect 3451 -2674 3485 -2640
rect 3519 -2674 3553 -2640
rect 3587 -2674 3621 -2640
rect 3655 -2674 3689 -2640
rect 3723 -2674 3757 -2640
rect 3791 -2674 3825 -2640
rect 3859 -2674 3893 -2640
rect 3927 -2674 3961 -2640
rect 3995 -2674 4029 -2640
rect 4063 -2674 4097 -2640
rect 4131 -2674 4247 -2640
<< psubdiffcont >>
rect -4131 2640 -4097 2674
rect -4063 2640 -4029 2674
rect -3995 2640 -3961 2674
rect -3927 2640 -3893 2674
rect -3859 2640 -3825 2674
rect -3791 2640 -3757 2674
rect -3723 2640 -3689 2674
rect -3655 2640 -3621 2674
rect -3587 2640 -3553 2674
rect -3519 2640 -3485 2674
rect -3451 2640 -3417 2674
rect -3383 2640 -3349 2674
rect -3315 2640 -3281 2674
rect -3247 2640 -3213 2674
rect -3179 2640 -3145 2674
rect -3111 2640 -3077 2674
rect -3043 2640 -3009 2674
rect -2975 2640 -2941 2674
rect -2907 2640 -2873 2674
rect -2839 2640 -2805 2674
rect -2771 2640 -2737 2674
rect -2703 2640 -2669 2674
rect -2635 2640 -2601 2674
rect -2567 2640 -2533 2674
rect -2499 2640 -2465 2674
rect -2431 2640 -2397 2674
rect -2363 2640 -2329 2674
rect -2295 2640 -2261 2674
rect -2227 2640 -2193 2674
rect -2159 2640 -2125 2674
rect -2091 2640 -2057 2674
rect -2023 2640 -1989 2674
rect -1955 2640 -1921 2674
rect -1887 2640 -1853 2674
rect -1819 2640 -1785 2674
rect -1751 2640 -1717 2674
rect -1683 2640 -1649 2674
rect -1615 2640 -1581 2674
rect -1547 2640 -1513 2674
rect -1479 2640 -1445 2674
rect -1411 2640 -1377 2674
rect -1343 2640 -1309 2674
rect -1275 2640 -1241 2674
rect -1207 2640 -1173 2674
rect -1139 2640 -1105 2674
rect -1071 2640 -1037 2674
rect -1003 2640 -969 2674
rect -935 2640 -901 2674
rect -867 2640 -833 2674
rect -799 2640 -765 2674
rect -731 2640 -697 2674
rect -663 2640 -629 2674
rect -595 2640 -561 2674
rect -527 2640 -493 2674
rect -459 2640 -425 2674
rect -391 2640 -357 2674
rect -323 2640 -289 2674
rect -255 2640 -221 2674
rect -187 2640 -153 2674
rect -119 2640 -85 2674
rect -51 2640 -17 2674
rect 17 2640 51 2674
rect 85 2640 119 2674
rect 153 2640 187 2674
rect 221 2640 255 2674
rect 289 2640 323 2674
rect 357 2640 391 2674
rect 425 2640 459 2674
rect 493 2640 527 2674
rect 561 2640 595 2674
rect 629 2640 663 2674
rect 697 2640 731 2674
rect 765 2640 799 2674
rect 833 2640 867 2674
rect 901 2640 935 2674
rect 969 2640 1003 2674
rect 1037 2640 1071 2674
rect 1105 2640 1139 2674
rect 1173 2640 1207 2674
rect 1241 2640 1275 2674
rect 1309 2640 1343 2674
rect 1377 2640 1411 2674
rect 1445 2640 1479 2674
rect 1513 2640 1547 2674
rect 1581 2640 1615 2674
rect 1649 2640 1683 2674
rect 1717 2640 1751 2674
rect 1785 2640 1819 2674
rect 1853 2640 1887 2674
rect 1921 2640 1955 2674
rect 1989 2640 2023 2674
rect 2057 2640 2091 2674
rect 2125 2640 2159 2674
rect 2193 2640 2227 2674
rect 2261 2640 2295 2674
rect 2329 2640 2363 2674
rect 2397 2640 2431 2674
rect 2465 2640 2499 2674
rect 2533 2640 2567 2674
rect 2601 2640 2635 2674
rect 2669 2640 2703 2674
rect 2737 2640 2771 2674
rect 2805 2640 2839 2674
rect 2873 2640 2907 2674
rect 2941 2640 2975 2674
rect 3009 2640 3043 2674
rect 3077 2640 3111 2674
rect 3145 2640 3179 2674
rect 3213 2640 3247 2674
rect 3281 2640 3315 2674
rect 3349 2640 3383 2674
rect 3417 2640 3451 2674
rect 3485 2640 3519 2674
rect 3553 2640 3587 2674
rect 3621 2640 3655 2674
rect 3689 2640 3723 2674
rect 3757 2640 3791 2674
rect 3825 2640 3859 2674
rect 3893 2640 3927 2674
rect 3961 2640 3995 2674
rect 4029 2640 4063 2674
rect 4097 2640 4131 2674
rect -4247 2533 -4213 2567
rect 4213 2533 4247 2567
rect -4247 2465 -4213 2499
rect -4247 2397 -4213 2431
rect -4247 2329 -4213 2363
rect -4247 2261 -4213 2295
rect -4247 2193 -4213 2227
rect -4247 2125 -4213 2159
rect -4247 2057 -4213 2091
rect -4247 1989 -4213 2023
rect -4247 1921 -4213 1955
rect -4247 1853 -4213 1887
rect -4247 1785 -4213 1819
rect -4247 1717 -4213 1751
rect -4247 1649 -4213 1683
rect -4247 1581 -4213 1615
rect -4247 1513 -4213 1547
rect -4247 1445 -4213 1479
rect -4247 1377 -4213 1411
rect -4247 1309 -4213 1343
rect -4247 1241 -4213 1275
rect -4247 1173 -4213 1207
rect -4247 1105 -4213 1139
rect -4247 1037 -4213 1071
rect -4247 969 -4213 1003
rect -4247 901 -4213 935
rect -4247 833 -4213 867
rect -4247 765 -4213 799
rect -4247 697 -4213 731
rect -4247 629 -4213 663
rect -4247 561 -4213 595
rect -4247 493 -4213 527
rect -4247 425 -4213 459
rect -4247 357 -4213 391
rect -4247 289 -4213 323
rect -4247 221 -4213 255
rect -4247 153 -4213 187
rect -4247 85 -4213 119
rect -4247 17 -4213 51
rect -4247 -51 -4213 -17
rect -4247 -119 -4213 -85
rect -4247 -187 -4213 -153
rect -4247 -255 -4213 -221
rect -4247 -323 -4213 -289
rect -4247 -391 -4213 -357
rect -4247 -459 -4213 -425
rect -4247 -527 -4213 -493
rect -4247 -595 -4213 -561
rect -4247 -663 -4213 -629
rect -4247 -731 -4213 -697
rect -4247 -799 -4213 -765
rect -4247 -867 -4213 -833
rect -4247 -935 -4213 -901
rect -4247 -1003 -4213 -969
rect -4247 -1071 -4213 -1037
rect -4247 -1139 -4213 -1105
rect -4247 -1207 -4213 -1173
rect -4247 -1275 -4213 -1241
rect -4247 -1343 -4213 -1309
rect -4247 -1411 -4213 -1377
rect -4247 -1479 -4213 -1445
rect -4247 -1547 -4213 -1513
rect -4247 -1615 -4213 -1581
rect -4247 -1683 -4213 -1649
rect -4247 -1751 -4213 -1717
rect -4247 -1819 -4213 -1785
rect -4247 -1887 -4213 -1853
rect -4247 -1955 -4213 -1921
rect -4247 -2023 -4213 -1989
rect -4247 -2091 -4213 -2057
rect -4247 -2159 -4213 -2125
rect -4247 -2227 -4213 -2193
rect -4247 -2295 -4213 -2261
rect -4247 -2363 -4213 -2329
rect -4247 -2431 -4213 -2397
rect -4247 -2499 -4213 -2465
rect 4213 2465 4247 2499
rect 4213 2397 4247 2431
rect 4213 2329 4247 2363
rect 4213 2261 4247 2295
rect 4213 2193 4247 2227
rect 4213 2125 4247 2159
rect 4213 2057 4247 2091
rect 4213 1989 4247 2023
rect 4213 1921 4247 1955
rect 4213 1853 4247 1887
rect 4213 1785 4247 1819
rect 4213 1717 4247 1751
rect 4213 1649 4247 1683
rect 4213 1581 4247 1615
rect 4213 1513 4247 1547
rect 4213 1445 4247 1479
rect 4213 1377 4247 1411
rect 4213 1309 4247 1343
rect 4213 1241 4247 1275
rect 4213 1173 4247 1207
rect 4213 1105 4247 1139
rect 4213 1037 4247 1071
rect 4213 969 4247 1003
rect 4213 901 4247 935
rect 4213 833 4247 867
rect 4213 765 4247 799
rect 4213 697 4247 731
rect 4213 629 4247 663
rect 4213 561 4247 595
rect 4213 493 4247 527
rect 4213 425 4247 459
rect 4213 357 4247 391
rect 4213 289 4247 323
rect 4213 221 4247 255
rect 4213 153 4247 187
rect 4213 85 4247 119
rect 4213 17 4247 51
rect 4213 -51 4247 -17
rect 4213 -119 4247 -85
rect 4213 -187 4247 -153
rect 4213 -255 4247 -221
rect 4213 -323 4247 -289
rect 4213 -391 4247 -357
rect 4213 -459 4247 -425
rect 4213 -527 4247 -493
rect 4213 -595 4247 -561
rect 4213 -663 4247 -629
rect 4213 -731 4247 -697
rect 4213 -799 4247 -765
rect 4213 -867 4247 -833
rect 4213 -935 4247 -901
rect 4213 -1003 4247 -969
rect 4213 -1071 4247 -1037
rect 4213 -1139 4247 -1105
rect 4213 -1207 4247 -1173
rect 4213 -1275 4247 -1241
rect 4213 -1343 4247 -1309
rect 4213 -1411 4247 -1377
rect 4213 -1479 4247 -1445
rect 4213 -1547 4247 -1513
rect 4213 -1615 4247 -1581
rect 4213 -1683 4247 -1649
rect 4213 -1751 4247 -1717
rect 4213 -1819 4247 -1785
rect 4213 -1887 4247 -1853
rect 4213 -1955 4247 -1921
rect 4213 -2023 4247 -1989
rect 4213 -2091 4247 -2057
rect 4213 -2159 4247 -2125
rect 4213 -2227 4247 -2193
rect 4213 -2295 4247 -2261
rect 4213 -2363 4247 -2329
rect 4213 -2431 4247 -2397
rect 4213 -2499 4247 -2465
rect -4247 -2567 -4213 -2533
rect 4213 -2567 4247 -2533
rect -4131 -2674 -4097 -2640
rect -4063 -2674 -4029 -2640
rect -3995 -2674 -3961 -2640
rect -3927 -2674 -3893 -2640
rect -3859 -2674 -3825 -2640
rect -3791 -2674 -3757 -2640
rect -3723 -2674 -3689 -2640
rect -3655 -2674 -3621 -2640
rect -3587 -2674 -3553 -2640
rect -3519 -2674 -3485 -2640
rect -3451 -2674 -3417 -2640
rect -3383 -2674 -3349 -2640
rect -3315 -2674 -3281 -2640
rect -3247 -2674 -3213 -2640
rect -3179 -2674 -3145 -2640
rect -3111 -2674 -3077 -2640
rect -3043 -2674 -3009 -2640
rect -2975 -2674 -2941 -2640
rect -2907 -2674 -2873 -2640
rect -2839 -2674 -2805 -2640
rect -2771 -2674 -2737 -2640
rect -2703 -2674 -2669 -2640
rect -2635 -2674 -2601 -2640
rect -2567 -2674 -2533 -2640
rect -2499 -2674 -2465 -2640
rect -2431 -2674 -2397 -2640
rect -2363 -2674 -2329 -2640
rect -2295 -2674 -2261 -2640
rect -2227 -2674 -2193 -2640
rect -2159 -2674 -2125 -2640
rect -2091 -2674 -2057 -2640
rect -2023 -2674 -1989 -2640
rect -1955 -2674 -1921 -2640
rect -1887 -2674 -1853 -2640
rect -1819 -2674 -1785 -2640
rect -1751 -2674 -1717 -2640
rect -1683 -2674 -1649 -2640
rect -1615 -2674 -1581 -2640
rect -1547 -2674 -1513 -2640
rect -1479 -2674 -1445 -2640
rect -1411 -2674 -1377 -2640
rect -1343 -2674 -1309 -2640
rect -1275 -2674 -1241 -2640
rect -1207 -2674 -1173 -2640
rect -1139 -2674 -1105 -2640
rect -1071 -2674 -1037 -2640
rect -1003 -2674 -969 -2640
rect -935 -2674 -901 -2640
rect -867 -2674 -833 -2640
rect -799 -2674 -765 -2640
rect -731 -2674 -697 -2640
rect -663 -2674 -629 -2640
rect -595 -2674 -561 -2640
rect -527 -2674 -493 -2640
rect -459 -2674 -425 -2640
rect -391 -2674 -357 -2640
rect -323 -2674 -289 -2640
rect -255 -2674 -221 -2640
rect -187 -2674 -153 -2640
rect -119 -2674 -85 -2640
rect -51 -2674 -17 -2640
rect 17 -2674 51 -2640
rect 85 -2674 119 -2640
rect 153 -2674 187 -2640
rect 221 -2674 255 -2640
rect 289 -2674 323 -2640
rect 357 -2674 391 -2640
rect 425 -2674 459 -2640
rect 493 -2674 527 -2640
rect 561 -2674 595 -2640
rect 629 -2674 663 -2640
rect 697 -2674 731 -2640
rect 765 -2674 799 -2640
rect 833 -2674 867 -2640
rect 901 -2674 935 -2640
rect 969 -2674 1003 -2640
rect 1037 -2674 1071 -2640
rect 1105 -2674 1139 -2640
rect 1173 -2674 1207 -2640
rect 1241 -2674 1275 -2640
rect 1309 -2674 1343 -2640
rect 1377 -2674 1411 -2640
rect 1445 -2674 1479 -2640
rect 1513 -2674 1547 -2640
rect 1581 -2674 1615 -2640
rect 1649 -2674 1683 -2640
rect 1717 -2674 1751 -2640
rect 1785 -2674 1819 -2640
rect 1853 -2674 1887 -2640
rect 1921 -2674 1955 -2640
rect 1989 -2674 2023 -2640
rect 2057 -2674 2091 -2640
rect 2125 -2674 2159 -2640
rect 2193 -2674 2227 -2640
rect 2261 -2674 2295 -2640
rect 2329 -2674 2363 -2640
rect 2397 -2674 2431 -2640
rect 2465 -2674 2499 -2640
rect 2533 -2674 2567 -2640
rect 2601 -2674 2635 -2640
rect 2669 -2674 2703 -2640
rect 2737 -2674 2771 -2640
rect 2805 -2674 2839 -2640
rect 2873 -2674 2907 -2640
rect 2941 -2674 2975 -2640
rect 3009 -2674 3043 -2640
rect 3077 -2674 3111 -2640
rect 3145 -2674 3179 -2640
rect 3213 -2674 3247 -2640
rect 3281 -2674 3315 -2640
rect 3349 -2674 3383 -2640
rect 3417 -2674 3451 -2640
rect 3485 -2674 3519 -2640
rect 3553 -2674 3587 -2640
rect 3621 -2674 3655 -2640
rect 3689 -2674 3723 -2640
rect 3757 -2674 3791 -2640
rect 3825 -2674 3859 -2640
rect 3893 -2674 3927 -2640
rect 3961 -2674 3995 -2640
rect 4029 -2674 4063 -2640
rect 4097 -2674 4131 -2640
<< poly >>
rect -4087 2572 -2087 2588
rect -4087 2538 -4056 2572
rect -4022 2538 -3988 2572
rect -3954 2538 -3920 2572
rect -3886 2538 -3852 2572
rect -3818 2538 -3784 2572
rect -3750 2538 -3716 2572
rect -3682 2538 -3648 2572
rect -3614 2538 -3580 2572
rect -3546 2538 -3512 2572
rect -3478 2538 -3444 2572
rect -3410 2538 -3376 2572
rect -3342 2538 -3308 2572
rect -3274 2538 -3240 2572
rect -3206 2538 -3172 2572
rect -3138 2538 -3104 2572
rect -3070 2538 -3036 2572
rect -3002 2538 -2968 2572
rect -2934 2538 -2900 2572
rect -2866 2538 -2832 2572
rect -2798 2538 -2764 2572
rect -2730 2538 -2696 2572
rect -2662 2538 -2628 2572
rect -2594 2538 -2560 2572
rect -2526 2538 -2492 2572
rect -2458 2538 -2424 2572
rect -2390 2538 -2356 2572
rect -2322 2538 -2288 2572
rect -2254 2538 -2220 2572
rect -2186 2538 -2152 2572
rect -2118 2538 -2087 2572
rect -4087 2500 -2087 2538
rect -2029 2572 -29 2588
rect -2029 2538 -1998 2572
rect -1964 2538 -1930 2572
rect -1896 2538 -1862 2572
rect -1828 2538 -1794 2572
rect -1760 2538 -1726 2572
rect -1692 2538 -1658 2572
rect -1624 2538 -1590 2572
rect -1556 2538 -1522 2572
rect -1488 2538 -1454 2572
rect -1420 2538 -1386 2572
rect -1352 2538 -1318 2572
rect -1284 2538 -1250 2572
rect -1216 2538 -1182 2572
rect -1148 2538 -1114 2572
rect -1080 2538 -1046 2572
rect -1012 2538 -978 2572
rect -944 2538 -910 2572
rect -876 2538 -842 2572
rect -808 2538 -774 2572
rect -740 2538 -706 2572
rect -672 2538 -638 2572
rect -604 2538 -570 2572
rect -536 2538 -502 2572
rect -468 2538 -434 2572
rect -400 2538 -366 2572
rect -332 2538 -298 2572
rect -264 2538 -230 2572
rect -196 2538 -162 2572
rect -128 2538 -94 2572
rect -60 2538 -29 2572
rect -2029 2500 -29 2538
rect 29 2572 2029 2588
rect 29 2538 60 2572
rect 94 2538 128 2572
rect 162 2538 196 2572
rect 230 2538 264 2572
rect 298 2538 332 2572
rect 366 2538 400 2572
rect 434 2538 468 2572
rect 502 2538 536 2572
rect 570 2538 604 2572
rect 638 2538 672 2572
rect 706 2538 740 2572
rect 774 2538 808 2572
rect 842 2538 876 2572
rect 910 2538 944 2572
rect 978 2538 1012 2572
rect 1046 2538 1080 2572
rect 1114 2538 1148 2572
rect 1182 2538 1216 2572
rect 1250 2538 1284 2572
rect 1318 2538 1352 2572
rect 1386 2538 1420 2572
rect 1454 2538 1488 2572
rect 1522 2538 1556 2572
rect 1590 2538 1624 2572
rect 1658 2538 1692 2572
rect 1726 2538 1760 2572
rect 1794 2538 1828 2572
rect 1862 2538 1896 2572
rect 1930 2538 1964 2572
rect 1998 2538 2029 2572
rect 29 2500 2029 2538
rect 2087 2572 4087 2588
rect 2087 2538 2118 2572
rect 2152 2538 2186 2572
rect 2220 2538 2254 2572
rect 2288 2538 2322 2572
rect 2356 2538 2390 2572
rect 2424 2538 2458 2572
rect 2492 2538 2526 2572
rect 2560 2538 2594 2572
rect 2628 2538 2662 2572
rect 2696 2538 2730 2572
rect 2764 2538 2798 2572
rect 2832 2538 2866 2572
rect 2900 2538 2934 2572
rect 2968 2538 3002 2572
rect 3036 2538 3070 2572
rect 3104 2538 3138 2572
rect 3172 2538 3206 2572
rect 3240 2538 3274 2572
rect 3308 2538 3342 2572
rect 3376 2538 3410 2572
rect 3444 2538 3478 2572
rect 3512 2538 3546 2572
rect 3580 2538 3614 2572
rect 3648 2538 3682 2572
rect 3716 2538 3750 2572
rect 3784 2538 3818 2572
rect 3852 2538 3886 2572
rect 3920 2538 3954 2572
rect 3988 2538 4022 2572
rect 4056 2538 4087 2572
rect 2087 2500 4087 2538
rect -4087 -2538 -2087 -2500
rect -4087 -2572 -4056 -2538
rect -4022 -2572 -3988 -2538
rect -3954 -2572 -3920 -2538
rect -3886 -2572 -3852 -2538
rect -3818 -2572 -3784 -2538
rect -3750 -2572 -3716 -2538
rect -3682 -2572 -3648 -2538
rect -3614 -2572 -3580 -2538
rect -3546 -2572 -3512 -2538
rect -3478 -2572 -3444 -2538
rect -3410 -2572 -3376 -2538
rect -3342 -2572 -3308 -2538
rect -3274 -2572 -3240 -2538
rect -3206 -2572 -3172 -2538
rect -3138 -2572 -3104 -2538
rect -3070 -2572 -3036 -2538
rect -3002 -2572 -2968 -2538
rect -2934 -2572 -2900 -2538
rect -2866 -2572 -2832 -2538
rect -2798 -2572 -2764 -2538
rect -2730 -2572 -2696 -2538
rect -2662 -2572 -2628 -2538
rect -2594 -2572 -2560 -2538
rect -2526 -2572 -2492 -2538
rect -2458 -2572 -2424 -2538
rect -2390 -2572 -2356 -2538
rect -2322 -2572 -2288 -2538
rect -2254 -2572 -2220 -2538
rect -2186 -2572 -2152 -2538
rect -2118 -2572 -2087 -2538
rect -4087 -2588 -2087 -2572
rect -2029 -2538 -29 -2500
rect -2029 -2572 -1998 -2538
rect -1964 -2572 -1930 -2538
rect -1896 -2572 -1862 -2538
rect -1828 -2572 -1794 -2538
rect -1760 -2572 -1726 -2538
rect -1692 -2572 -1658 -2538
rect -1624 -2572 -1590 -2538
rect -1556 -2572 -1522 -2538
rect -1488 -2572 -1454 -2538
rect -1420 -2572 -1386 -2538
rect -1352 -2572 -1318 -2538
rect -1284 -2572 -1250 -2538
rect -1216 -2572 -1182 -2538
rect -1148 -2572 -1114 -2538
rect -1080 -2572 -1046 -2538
rect -1012 -2572 -978 -2538
rect -944 -2572 -910 -2538
rect -876 -2572 -842 -2538
rect -808 -2572 -774 -2538
rect -740 -2572 -706 -2538
rect -672 -2572 -638 -2538
rect -604 -2572 -570 -2538
rect -536 -2572 -502 -2538
rect -468 -2572 -434 -2538
rect -400 -2572 -366 -2538
rect -332 -2572 -298 -2538
rect -264 -2572 -230 -2538
rect -196 -2572 -162 -2538
rect -128 -2572 -94 -2538
rect -60 -2572 -29 -2538
rect -2029 -2588 -29 -2572
rect 29 -2538 2029 -2500
rect 29 -2572 60 -2538
rect 94 -2572 128 -2538
rect 162 -2572 196 -2538
rect 230 -2572 264 -2538
rect 298 -2572 332 -2538
rect 366 -2572 400 -2538
rect 434 -2572 468 -2538
rect 502 -2572 536 -2538
rect 570 -2572 604 -2538
rect 638 -2572 672 -2538
rect 706 -2572 740 -2538
rect 774 -2572 808 -2538
rect 842 -2572 876 -2538
rect 910 -2572 944 -2538
rect 978 -2572 1012 -2538
rect 1046 -2572 1080 -2538
rect 1114 -2572 1148 -2538
rect 1182 -2572 1216 -2538
rect 1250 -2572 1284 -2538
rect 1318 -2572 1352 -2538
rect 1386 -2572 1420 -2538
rect 1454 -2572 1488 -2538
rect 1522 -2572 1556 -2538
rect 1590 -2572 1624 -2538
rect 1658 -2572 1692 -2538
rect 1726 -2572 1760 -2538
rect 1794 -2572 1828 -2538
rect 1862 -2572 1896 -2538
rect 1930 -2572 1964 -2538
rect 1998 -2572 2029 -2538
rect 29 -2588 2029 -2572
rect 2087 -2538 4087 -2500
rect 2087 -2572 2118 -2538
rect 2152 -2572 2186 -2538
rect 2220 -2572 2254 -2538
rect 2288 -2572 2322 -2538
rect 2356 -2572 2390 -2538
rect 2424 -2572 2458 -2538
rect 2492 -2572 2526 -2538
rect 2560 -2572 2594 -2538
rect 2628 -2572 2662 -2538
rect 2696 -2572 2730 -2538
rect 2764 -2572 2798 -2538
rect 2832 -2572 2866 -2538
rect 2900 -2572 2934 -2538
rect 2968 -2572 3002 -2538
rect 3036 -2572 3070 -2538
rect 3104 -2572 3138 -2538
rect 3172 -2572 3206 -2538
rect 3240 -2572 3274 -2538
rect 3308 -2572 3342 -2538
rect 3376 -2572 3410 -2538
rect 3444 -2572 3478 -2538
rect 3512 -2572 3546 -2538
rect 3580 -2572 3614 -2538
rect 3648 -2572 3682 -2538
rect 3716 -2572 3750 -2538
rect 3784 -2572 3818 -2538
rect 3852 -2572 3886 -2538
rect 3920 -2572 3954 -2538
rect 3988 -2572 4022 -2538
rect 4056 -2572 4087 -2538
rect 2087 -2588 4087 -2572
<< polycont >>
rect -4056 2538 -4022 2572
rect -3988 2538 -3954 2572
rect -3920 2538 -3886 2572
rect -3852 2538 -3818 2572
rect -3784 2538 -3750 2572
rect -3716 2538 -3682 2572
rect -3648 2538 -3614 2572
rect -3580 2538 -3546 2572
rect -3512 2538 -3478 2572
rect -3444 2538 -3410 2572
rect -3376 2538 -3342 2572
rect -3308 2538 -3274 2572
rect -3240 2538 -3206 2572
rect -3172 2538 -3138 2572
rect -3104 2538 -3070 2572
rect -3036 2538 -3002 2572
rect -2968 2538 -2934 2572
rect -2900 2538 -2866 2572
rect -2832 2538 -2798 2572
rect -2764 2538 -2730 2572
rect -2696 2538 -2662 2572
rect -2628 2538 -2594 2572
rect -2560 2538 -2526 2572
rect -2492 2538 -2458 2572
rect -2424 2538 -2390 2572
rect -2356 2538 -2322 2572
rect -2288 2538 -2254 2572
rect -2220 2538 -2186 2572
rect -2152 2538 -2118 2572
rect -1998 2538 -1964 2572
rect -1930 2538 -1896 2572
rect -1862 2538 -1828 2572
rect -1794 2538 -1760 2572
rect -1726 2538 -1692 2572
rect -1658 2538 -1624 2572
rect -1590 2538 -1556 2572
rect -1522 2538 -1488 2572
rect -1454 2538 -1420 2572
rect -1386 2538 -1352 2572
rect -1318 2538 -1284 2572
rect -1250 2538 -1216 2572
rect -1182 2538 -1148 2572
rect -1114 2538 -1080 2572
rect -1046 2538 -1012 2572
rect -978 2538 -944 2572
rect -910 2538 -876 2572
rect -842 2538 -808 2572
rect -774 2538 -740 2572
rect -706 2538 -672 2572
rect -638 2538 -604 2572
rect -570 2538 -536 2572
rect -502 2538 -468 2572
rect -434 2538 -400 2572
rect -366 2538 -332 2572
rect -298 2538 -264 2572
rect -230 2538 -196 2572
rect -162 2538 -128 2572
rect -94 2538 -60 2572
rect 60 2538 94 2572
rect 128 2538 162 2572
rect 196 2538 230 2572
rect 264 2538 298 2572
rect 332 2538 366 2572
rect 400 2538 434 2572
rect 468 2538 502 2572
rect 536 2538 570 2572
rect 604 2538 638 2572
rect 672 2538 706 2572
rect 740 2538 774 2572
rect 808 2538 842 2572
rect 876 2538 910 2572
rect 944 2538 978 2572
rect 1012 2538 1046 2572
rect 1080 2538 1114 2572
rect 1148 2538 1182 2572
rect 1216 2538 1250 2572
rect 1284 2538 1318 2572
rect 1352 2538 1386 2572
rect 1420 2538 1454 2572
rect 1488 2538 1522 2572
rect 1556 2538 1590 2572
rect 1624 2538 1658 2572
rect 1692 2538 1726 2572
rect 1760 2538 1794 2572
rect 1828 2538 1862 2572
rect 1896 2538 1930 2572
rect 1964 2538 1998 2572
rect 2118 2538 2152 2572
rect 2186 2538 2220 2572
rect 2254 2538 2288 2572
rect 2322 2538 2356 2572
rect 2390 2538 2424 2572
rect 2458 2538 2492 2572
rect 2526 2538 2560 2572
rect 2594 2538 2628 2572
rect 2662 2538 2696 2572
rect 2730 2538 2764 2572
rect 2798 2538 2832 2572
rect 2866 2538 2900 2572
rect 2934 2538 2968 2572
rect 3002 2538 3036 2572
rect 3070 2538 3104 2572
rect 3138 2538 3172 2572
rect 3206 2538 3240 2572
rect 3274 2538 3308 2572
rect 3342 2538 3376 2572
rect 3410 2538 3444 2572
rect 3478 2538 3512 2572
rect 3546 2538 3580 2572
rect 3614 2538 3648 2572
rect 3682 2538 3716 2572
rect 3750 2538 3784 2572
rect 3818 2538 3852 2572
rect 3886 2538 3920 2572
rect 3954 2538 3988 2572
rect 4022 2538 4056 2572
rect -4056 -2572 -4022 -2538
rect -3988 -2572 -3954 -2538
rect -3920 -2572 -3886 -2538
rect -3852 -2572 -3818 -2538
rect -3784 -2572 -3750 -2538
rect -3716 -2572 -3682 -2538
rect -3648 -2572 -3614 -2538
rect -3580 -2572 -3546 -2538
rect -3512 -2572 -3478 -2538
rect -3444 -2572 -3410 -2538
rect -3376 -2572 -3342 -2538
rect -3308 -2572 -3274 -2538
rect -3240 -2572 -3206 -2538
rect -3172 -2572 -3138 -2538
rect -3104 -2572 -3070 -2538
rect -3036 -2572 -3002 -2538
rect -2968 -2572 -2934 -2538
rect -2900 -2572 -2866 -2538
rect -2832 -2572 -2798 -2538
rect -2764 -2572 -2730 -2538
rect -2696 -2572 -2662 -2538
rect -2628 -2572 -2594 -2538
rect -2560 -2572 -2526 -2538
rect -2492 -2572 -2458 -2538
rect -2424 -2572 -2390 -2538
rect -2356 -2572 -2322 -2538
rect -2288 -2572 -2254 -2538
rect -2220 -2572 -2186 -2538
rect -2152 -2572 -2118 -2538
rect -1998 -2572 -1964 -2538
rect -1930 -2572 -1896 -2538
rect -1862 -2572 -1828 -2538
rect -1794 -2572 -1760 -2538
rect -1726 -2572 -1692 -2538
rect -1658 -2572 -1624 -2538
rect -1590 -2572 -1556 -2538
rect -1522 -2572 -1488 -2538
rect -1454 -2572 -1420 -2538
rect -1386 -2572 -1352 -2538
rect -1318 -2572 -1284 -2538
rect -1250 -2572 -1216 -2538
rect -1182 -2572 -1148 -2538
rect -1114 -2572 -1080 -2538
rect -1046 -2572 -1012 -2538
rect -978 -2572 -944 -2538
rect -910 -2572 -876 -2538
rect -842 -2572 -808 -2538
rect -774 -2572 -740 -2538
rect -706 -2572 -672 -2538
rect -638 -2572 -604 -2538
rect -570 -2572 -536 -2538
rect -502 -2572 -468 -2538
rect -434 -2572 -400 -2538
rect -366 -2572 -332 -2538
rect -298 -2572 -264 -2538
rect -230 -2572 -196 -2538
rect -162 -2572 -128 -2538
rect -94 -2572 -60 -2538
rect 60 -2572 94 -2538
rect 128 -2572 162 -2538
rect 196 -2572 230 -2538
rect 264 -2572 298 -2538
rect 332 -2572 366 -2538
rect 400 -2572 434 -2538
rect 468 -2572 502 -2538
rect 536 -2572 570 -2538
rect 604 -2572 638 -2538
rect 672 -2572 706 -2538
rect 740 -2572 774 -2538
rect 808 -2572 842 -2538
rect 876 -2572 910 -2538
rect 944 -2572 978 -2538
rect 1012 -2572 1046 -2538
rect 1080 -2572 1114 -2538
rect 1148 -2572 1182 -2538
rect 1216 -2572 1250 -2538
rect 1284 -2572 1318 -2538
rect 1352 -2572 1386 -2538
rect 1420 -2572 1454 -2538
rect 1488 -2572 1522 -2538
rect 1556 -2572 1590 -2538
rect 1624 -2572 1658 -2538
rect 1692 -2572 1726 -2538
rect 1760 -2572 1794 -2538
rect 1828 -2572 1862 -2538
rect 1896 -2572 1930 -2538
rect 1964 -2572 1998 -2538
rect 2118 -2572 2152 -2538
rect 2186 -2572 2220 -2538
rect 2254 -2572 2288 -2538
rect 2322 -2572 2356 -2538
rect 2390 -2572 2424 -2538
rect 2458 -2572 2492 -2538
rect 2526 -2572 2560 -2538
rect 2594 -2572 2628 -2538
rect 2662 -2572 2696 -2538
rect 2730 -2572 2764 -2538
rect 2798 -2572 2832 -2538
rect 2866 -2572 2900 -2538
rect 2934 -2572 2968 -2538
rect 3002 -2572 3036 -2538
rect 3070 -2572 3104 -2538
rect 3138 -2572 3172 -2538
rect 3206 -2572 3240 -2538
rect 3274 -2572 3308 -2538
rect 3342 -2572 3376 -2538
rect 3410 -2572 3444 -2538
rect 3478 -2572 3512 -2538
rect 3546 -2572 3580 -2538
rect 3614 -2572 3648 -2538
rect 3682 -2572 3716 -2538
rect 3750 -2572 3784 -2538
rect 3818 -2572 3852 -2538
rect 3886 -2572 3920 -2538
rect 3954 -2572 3988 -2538
rect 4022 -2572 4056 -2538
<< locali >>
rect -4247 2640 -4131 2674
rect -4097 2640 -4063 2674
rect -4029 2640 -3995 2674
rect -3961 2640 -3927 2674
rect -3893 2640 -3859 2674
rect -3825 2640 -3791 2674
rect -3757 2640 -3723 2674
rect -3689 2640 -3655 2674
rect -3621 2640 -3587 2674
rect -3553 2640 -3519 2674
rect -3485 2640 -3451 2674
rect -3417 2640 -3383 2674
rect -3349 2640 -3315 2674
rect -3281 2640 -3247 2674
rect -3213 2640 -3179 2674
rect -3145 2640 -3111 2674
rect -3077 2640 -3043 2674
rect -3009 2640 -2975 2674
rect -2941 2640 -2907 2674
rect -2873 2640 -2839 2674
rect -2805 2640 -2771 2674
rect -2737 2640 -2703 2674
rect -2669 2640 -2635 2674
rect -2601 2640 -2567 2674
rect -2533 2640 -2499 2674
rect -2465 2640 -2431 2674
rect -2397 2640 -2363 2674
rect -2329 2640 -2295 2674
rect -2261 2640 -2227 2674
rect -2193 2640 -2159 2674
rect -2125 2640 -2091 2674
rect -2057 2640 -2023 2674
rect -1989 2640 -1955 2674
rect -1921 2640 -1887 2674
rect -1853 2640 -1819 2674
rect -1785 2640 -1751 2674
rect -1717 2640 -1683 2674
rect -1649 2640 -1615 2674
rect -1581 2640 -1547 2674
rect -1513 2640 -1479 2674
rect -1445 2640 -1411 2674
rect -1377 2640 -1343 2674
rect -1309 2640 -1275 2674
rect -1241 2640 -1207 2674
rect -1173 2640 -1139 2674
rect -1105 2640 -1071 2674
rect -1037 2640 -1003 2674
rect -969 2640 -935 2674
rect -901 2640 -867 2674
rect -833 2640 -799 2674
rect -765 2640 -731 2674
rect -697 2640 -663 2674
rect -629 2640 -595 2674
rect -561 2640 -527 2674
rect -493 2640 -459 2674
rect -425 2640 -391 2674
rect -357 2640 -323 2674
rect -289 2640 -255 2674
rect -221 2640 -187 2674
rect -153 2640 -119 2674
rect -85 2640 -51 2674
rect -17 2640 17 2674
rect 51 2640 85 2674
rect 119 2640 153 2674
rect 187 2640 221 2674
rect 255 2640 289 2674
rect 323 2640 357 2674
rect 391 2640 425 2674
rect 459 2640 493 2674
rect 527 2640 561 2674
rect 595 2640 629 2674
rect 663 2640 697 2674
rect 731 2640 765 2674
rect 799 2640 833 2674
rect 867 2640 901 2674
rect 935 2640 969 2674
rect 1003 2640 1037 2674
rect 1071 2640 1105 2674
rect 1139 2640 1173 2674
rect 1207 2640 1241 2674
rect 1275 2640 1309 2674
rect 1343 2640 1377 2674
rect 1411 2640 1445 2674
rect 1479 2640 1513 2674
rect 1547 2640 1581 2674
rect 1615 2640 1649 2674
rect 1683 2640 1717 2674
rect 1751 2640 1785 2674
rect 1819 2640 1853 2674
rect 1887 2640 1921 2674
rect 1955 2640 1989 2674
rect 2023 2640 2057 2674
rect 2091 2640 2125 2674
rect 2159 2640 2193 2674
rect 2227 2640 2261 2674
rect 2295 2640 2329 2674
rect 2363 2640 2397 2674
rect 2431 2640 2465 2674
rect 2499 2640 2533 2674
rect 2567 2640 2601 2674
rect 2635 2640 2669 2674
rect 2703 2640 2737 2674
rect 2771 2640 2805 2674
rect 2839 2640 2873 2674
rect 2907 2640 2941 2674
rect 2975 2640 3009 2674
rect 3043 2640 3077 2674
rect 3111 2640 3145 2674
rect 3179 2640 3213 2674
rect 3247 2640 3281 2674
rect 3315 2640 3349 2674
rect 3383 2640 3417 2674
rect 3451 2640 3485 2674
rect 3519 2640 3553 2674
rect 3587 2640 3621 2674
rect 3655 2640 3689 2674
rect 3723 2640 3757 2674
rect 3791 2640 3825 2674
rect 3859 2640 3893 2674
rect 3927 2640 3961 2674
rect 3995 2640 4029 2674
rect 4063 2640 4097 2674
rect 4131 2640 4247 2674
rect -4247 2567 -4213 2640
rect -4087 2538 -4056 2572
rect -4006 2538 -3988 2572
rect -3934 2538 -3920 2572
rect -3862 2538 -3852 2572
rect -3790 2538 -3784 2572
rect -3718 2538 -3716 2572
rect -3682 2538 -3680 2572
rect -3614 2538 -3608 2572
rect -3546 2538 -3536 2572
rect -3478 2538 -3464 2572
rect -3410 2538 -3392 2572
rect -3342 2538 -3320 2572
rect -3274 2538 -3248 2572
rect -3206 2538 -3176 2572
rect -3138 2538 -3104 2572
rect -3070 2538 -3036 2572
rect -2998 2538 -2968 2572
rect -2926 2538 -2900 2572
rect -2854 2538 -2832 2572
rect -2782 2538 -2764 2572
rect -2710 2538 -2696 2572
rect -2638 2538 -2628 2572
rect -2566 2538 -2560 2572
rect -2494 2538 -2492 2572
rect -2458 2538 -2456 2572
rect -2390 2538 -2384 2572
rect -2322 2538 -2312 2572
rect -2254 2538 -2240 2572
rect -2186 2538 -2168 2572
rect -2118 2538 -2087 2572
rect -2029 2538 -1998 2572
rect -1948 2538 -1930 2572
rect -1876 2538 -1862 2572
rect -1804 2538 -1794 2572
rect -1732 2538 -1726 2572
rect -1660 2538 -1658 2572
rect -1624 2538 -1622 2572
rect -1556 2538 -1550 2572
rect -1488 2538 -1478 2572
rect -1420 2538 -1406 2572
rect -1352 2538 -1334 2572
rect -1284 2538 -1262 2572
rect -1216 2538 -1190 2572
rect -1148 2538 -1118 2572
rect -1080 2538 -1046 2572
rect -1012 2538 -978 2572
rect -940 2538 -910 2572
rect -868 2538 -842 2572
rect -796 2538 -774 2572
rect -724 2538 -706 2572
rect -652 2538 -638 2572
rect -580 2538 -570 2572
rect -508 2538 -502 2572
rect -436 2538 -434 2572
rect -400 2538 -398 2572
rect -332 2538 -326 2572
rect -264 2538 -254 2572
rect -196 2538 -182 2572
rect -128 2538 -110 2572
rect -60 2538 -29 2572
rect 29 2538 60 2572
rect 110 2538 128 2572
rect 182 2538 196 2572
rect 254 2538 264 2572
rect 326 2538 332 2572
rect 398 2538 400 2572
rect 434 2538 436 2572
rect 502 2538 508 2572
rect 570 2538 580 2572
rect 638 2538 652 2572
rect 706 2538 724 2572
rect 774 2538 796 2572
rect 842 2538 868 2572
rect 910 2538 940 2572
rect 978 2538 1012 2572
rect 1046 2538 1080 2572
rect 1118 2538 1148 2572
rect 1190 2538 1216 2572
rect 1262 2538 1284 2572
rect 1334 2538 1352 2572
rect 1406 2538 1420 2572
rect 1478 2538 1488 2572
rect 1550 2538 1556 2572
rect 1622 2538 1624 2572
rect 1658 2538 1660 2572
rect 1726 2538 1732 2572
rect 1794 2538 1804 2572
rect 1862 2538 1876 2572
rect 1930 2538 1948 2572
rect 1998 2538 2029 2572
rect 2087 2538 2118 2572
rect 2168 2538 2186 2572
rect 2240 2538 2254 2572
rect 2312 2538 2322 2572
rect 2384 2538 2390 2572
rect 2456 2538 2458 2572
rect 2492 2538 2494 2572
rect 2560 2538 2566 2572
rect 2628 2538 2638 2572
rect 2696 2538 2710 2572
rect 2764 2538 2782 2572
rect 2832 2538 2854 2572
rect 2900 2538 2926 2572
rect 2968 2538 2998 2572
rect 3036 2538 3070 2572
rect 3104 2538 3138 2572
rect 3176 2538 3206 2572
rect 3248 2538 3274 2572
rect 3320 2538 3342 2572
rect 3392 2538 3410 2572
rect 3464 2538 3478 2572
rect 3536 2538 3546 2572
rect 3608 2538 3614 2572
rect 3680 2538 3682 2572
rect 3716 2538 3718 2572
rect 3784 2538 3790 2572
rect 3852 2538 3862 2572
rect 3920 2538 3934 2572
rect 3988 2538 4006 2572
rect 4056 2538 4087 2572
rect 4213 2567 4247 2640
rect -4247 2499 -4213 2533
rect -4247 2431 -4213 2465
rect -4247 2363 -4213 2397
rect -4247 2295 -4213 2329
rect -4247 2227 -4213 2261
rect -4247 2159 -4213 2193
rect -4247 2091 -4213 2125
rect -4247 2023 -4213 2057
rect -4247 1955 -4213 1989
rect -4247 1887 -4213 1921
rect -4247 1819 -4213 1853
rect -4247 1751 -4213 1785
rect -4247 1683 -4213 1717
rect -4247 1615 -4213 1649
rect -4247 1547 -4213 1581
rect -4247 1479 -4213 1513
rect -4247 1411 -4213 1445
rect -4247 1343 -4213 1377
rect -4247 1275 -4213 1309
rect -4247 1207 -4213 1241
rect -4247 1139 -4213 1173
rect -4247 1071 -4213 1105
rect -4247 1003 -4213 1037
rect -4247 935 -4213 969
rect -4247 867 -4213 901
rect -4247 799 -4213 833
rect -4247 731 -4213 765
rect -4247 663 -4213 697
rect -4247 595 -4213 629
rect -4247 527 -4213 561
rect -4247 459 -4213 493
rect -4247 391 -4213 425
rect -4247 323 -4213 357
rect -4247 255 -4213 289
rect -4247 187 -4213 221
rect -4247 119 -4213 153
rect -4247 51 -4213 85
rect -4247 -17 -4213 17
rect -4247 -85 -4213 -51
rect -4247 -153 -4213 -119
rect -4247 -221 -4213 -187
rect -4247 -289 -4213 -255
rect -4247 -357 -4213 -323
rect -4247 -425 -4213 -391
rect -4247 -493 -4213 -459
rect -4247 -561 -4213 -527
rect -4247 -629 -4213 -595
rect -4247 -697 -4213 -663
rect -4247 -765 -4213 -731
rect -4247 -833 -4213 -799
rect -4247 -901 -4213 -867
rect -4247 -969 -4213 -935
rect -4247 -1037 -4213 -1003
rect -4247 -1105 -4213 -1071
rect -4247 -1173 -4213 -1139
rect -4247 -1241 -4213 -1207
rect -4247 -1309 -4213 -1275
rect -4247 -1377 -4213 -1343
rect -4247 -1445 -4213 -1411
rect -4247 -1513 -4213 -1479
rect -4247 -1581 -4213 -1547
rect -4247 -1649 -4213 -1615
rect -4247 -1717 -4213 -1683
rect -4247 -1785 -4213 -1751
rect -4247 -1853 -4213 -1819
rect -4247 -1921 -4213 -1887
rect -4247 -1989 -4213 -1955
rect -4247 -2057 -4213 -2023
rect -4247 -2125 -4213 -2091
rect -4247 -2193 -4213 -2159
rect -4247 -2261 -4213 -2227
rect -4247 -2329 -4213 -2295
rect -4247 -2397 -4213 -2363
rect -4247 -2465 -4213 -2431
rect -4247 -2533 -4213 -2499
rect -4133 2465 -4099 2504
rect -4133 2397 -4099 2431
rect -4133 2329 -4099 2359
rect -4133 2261 -4099 2287
rect -4133 2193 -4099 2215
rect -4133 2125 -4099 2143
rect -4133 2057 -4099 2071
rect -4133 1989 -4099 1999
rect -4133 1921 -4099 1927
rect -4133 1853 -4099 1855
rect -4133 1817 -4099 1819
rect -4133 1745 -4099 1751
rect -4133 1673 -4099 1683
rect -4133 1601 -4099 1615
rect -4133 1529 -4099 1547
rect -4133 1457 -4099 1479
rect -4133 1385 -4099 1411
rect -4133 1313 -4099 1343
rect -4133 1241 -4099 1275
rect -4133 1173 -4099 1207
rect -4133 1105 -4099 1135
rect -4133 1037 -4099 1063
rect -4133 969 -4099 991
rect -4133 901 -4099 919
rect -4133 833 -4099 847
rect -4133 765 -4099 775
rect -4133 697 -4099 703
rect -4133 629 -4099 631
rect -4133 593 -4099 595
rect -4133 521 -4099 527
rect -4133 449 -4099 459
rect -4133 377 -4099 391
rect -4133 305 -4099 323
rect -4133 233 -4099 255
rect -4133 161 -4099 187
rect -4133 89 -4099 119
rect -4133 17 -4099 51
rect -4133 -51 -4099 -17
rect -4133 -119 -4099 -89
rect -4133 -187 -4099 -161
rect -4133 -255 -4099 -233
rect -4133 -323 -4099 -305
rect -4133 -391 -4099 -377
rect -4133 -459 -4099 -449
rect -4133 -527 -4099 -521
rect -4133 -595 -4099 -593
rect -4133 -631 -4099 -629
rect -4133 -703 -4099 -697
rect -4133 -775 -4099 -765
rect -4133 -847 -4099 -833
rect -4133 -919 -4099 -901
rect -4133 -991 -4099 -969
rect -4133 -1063 -4099 -1037
rect -4133 -1135 -4099 -1105
rect -4133 -1207 -4099 -1173
rect -4133 -1275 -4099 -1241
rect -4133 -1343 -4099 -1313
rect -4133 -1411 -4099 -1385
rect -4133 -1479 -4099 -1457
rect -4133 -1547 -4099 -1529
rect -4133 -1615 -4099 -1601
rect -4133 -1683 -4099 -1673
rect -4133 -1751 -4099 -1745
rect -4133 -1819 -4099 -1817
rect -4133 -1855 -4099 -1853
rect -4133 -1927 -4099 -1921
rect -4133 -1999 -4099 -1989
rect -4133 -2071 -4099 -2057
rect -4133 -2143 -4099 -2125
rect -4133 -2215 -4099 -2193
rect -4133 -2287 -4099 -2261
rect -4133 -2359 -4099 -2329
rect -4133 -2431 -4099 -2397
rect -4133 -2504 -4099 -2465
rect -2075 2465 -2041 2504
rect -2075 2397 -2041 2431
rect -2075 2329 -2041 2359
rect -2075 2261 -2041 2287
rect -2075 2193 -2041 2215
rect -2075 2125 -2041 2143
rect -2075 2057 -2041 2071
rect -2075 1989 -2041 1999
rect -2075 1921 -2041 1927
rect -2075 1853 -2041 1855
rect -2075 1817 -2041 1819
rect -2075 1745 -2041 1751
rect -2075 1673 -2041 1683
rect -2075 1601 -2041 1615
rect -2075 1529 -2041 1547
rect -2075 1457 -2041 1479
rect -2075 1385 -2041 1411
rect -2075 1313 -2041 1343
rect -2075 1241 -2041 1275
rect -2075 1173 -2041 1207
rect -2075 1105 -2041 1135
rect -2075 1037 -2041 1063
rect -2075 969 -2041 991
rect -2075 901 -2041 919
rect -2075 833 -2041 847
rect -2075 765 -2041 775
rect -2075 697 -2041 703
rect -2075 629 -2041 631
rect -2075 593 -2041 595
rect -2075 521 -2041 527
rect -2075 449 -2041 459
rect -2075 377 -2041 391
rect -2075 305 -2041 323
rect -2075 233 -2041 255
rect -2075 161 -2041 187
rect -2075 89 -2041 119
rect -2075 17 -2041 51
rect -2075 -51 -2041 -17
rect -2075 -119 -2041 -89
rect -2075 -187 -2041 -161
rect -2075 -255 -2041 -233
rect -2075 -323 -2041 -305
rect -2075 -391 -2041 -377
rect -2075 -459 -2041 -449
rect -2075 -527 -2041 -521
rect -2075 -595 -2041 -593
rect -2075 -631 -2041 -629
rect -2075 -703 -2041 -697
rect -2075 -775 -2041 -765
rect -2075 -847 -2041 -833
rect -2075 -919 -2041 -901
rect -2075 -991 -2041 -969
rect -2075 -1063 -2041 -1037
rect -2075 -1135 -2041 -1105
rect -2075 -1207 -2041 -1173
rect -2075 -1275 -2041 -1241
rect -2075 -1343 -2041 -1313
rect -2075 -1411 -2041 -1385
rect -2075 -1479 -2041 -1457
rect -2075 -1547 -2041 -1529
rect -2075 -1615 -2041 -1601
rect -2075 -1683 -2041 -1673
rect -2075 -1751 -2041 -1745
rect -2075 -1819 -2041 -1817
rect -2075 -1855 -2041 -1853
rect -2075 -1927 -2041 -1921
rect -2075 -1999 -2041 -1989
rect -2075 -2071 -2041 -2057
rect -2075 -2143 -2041 -2125
rect -2075 -2215 -2041 -2193
rect -2075 -2287 -2041 -2261
rect -2075 -2359 -2041 -2329
rect -2075 -2431 -2041 -2397
rect -2075 -2504 -2041 -2465
rect -17 2465 17 2504
rect -17 2397 17 2431
rect -17 2329 17 2359
rect -17 2261 17 2287
rect -17 2193 17 2215
rect -17 2125 17 2143
rect -17 2057 17 2071
rect -17 1989 17 1999
rect -17 1921 17 1927
rect -17 1853 17 1855
rect -17 1817 17 1819
rect -17 1745 17 1751
rect -17 1673 17 1683
rect -17 1601 17 1615
rect -17 1529 17 1547
rect -17 1457 17 1479
rect -17 1385 17 1411
rect -17 1313 17 1343
rect -17 1241 17 1275
rect -17 1173 17 1207
rect -17 1105 17 1135
rect -17 1037 17 1063
rect -17 969 17 991
rect -17 901 17 919
rect -17 833 17 847
rect -17 765 17 775
rect -17 697 17 703
rect -17 629 17 631
rect -17 593 17 595
rect -17 521 17 527
rect -17 449 17 459
rect -17 377 17 391
rect -17 305 17 323
rect -17 233 17 255
rect -17 161 17 187
rect -17 89 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -89
rect -17 -187 17 -161
rect -17 -255 17 -233
rect -17 -323 17 -305
rect -17 -391 17 -377
rect -17 -459 17 -449
rect -17 -527 17 -521
rect -17 -595 17 -593
rect -17 -631 17 -629
rect -17 -703 17 -697
rect -17 -775 17 -765
rect -17 -847 17 -833
rect -17 -919 17 -901
rect -17 -991 17 -969
rect -17 -1063 17 -1037
rect -17 -1135 17 -1105
rect -17 -1207 17 -1173
rect -17 -1275 17 -1241
rect -17 -1343 17 -1313
rect -17 -1411 17 -1385
rect -17 -1479 17 -1457
rect -17 -1547 17 -1529
rect -17 -1615 17 -1601
rect -17 -1683 17 -1673
rect -17 -1751 17 -1745
rect -17 -1819 17 -1817
rect -17 -1855 17 -1853
rect -17 -1927 17 -1921
rect -17 -1999 17 -1989
rect -17 -2071 17 -2057
rect -17 -2143 17 -2125
rect -17 -2215 17 -2193
rect -17 -2287 17 -2261
rect -17 -2359 17 -2329
rect -17 -2431 17 -2397
rect -17 -2504 17 -2465
rect 2041 2465 2075 2504
rect 2041 2397 2075 2431
rect 2041 2329 2075 2359
rect 2041 2261 2075 2287
rect 2041 2193 2075 2215
rect 2041 2125 2075 2143
rect 2041 2057 2075 2071
rect 2041 1989 2075 1999
rect 2041 1921 2075 1927
rect 2041 1853 2075 1855
rect 2041 1817 2075 1819
rect 2041 1745 2075 1751
rect 2041 1673 2075 1683
rect 2041 1601 2075 1615
rect 2041 1529 2075 1547
rect 2041 1457 2075 1479
rect 2041 1385 2075 1411
rect 2041 1313 2075 1343
rect 2041 1241 2075 1275
rect 2041 1173 2075 1207
rect 2041 1105 2075 1135
rect 2041 1037 2075 1063
rect 2041 969 2075 991
rect 2041 901 2075 919
rect 2041 833 2075 847
rect 2041 765 2075 775
rect 2041 697 2075 703
rect 2041 629 2075 631
rect 2041 593 2075 595
rect 2041 521 2075 527
rect 2041 449 2075 459
rect 2041 377 2075 391
rect 2041 305 2075 323
rect 2041 233 2075 255
rect 2041 161 2075 187
rect 2041 89 2075 119
rect 2041 17 2075 51
rect 2041 -51 2075 -17
rect 2041 -119 2075 -89
rect 2041 -187 2075 -161
rect 2041 -255 2075 -233
rect 2041 -323 2075 -305
rect 2041 -391 2075 -377
rect 2041 -459 2075 -449
rect 2041 -527 2075 -521
rect 2041 -595 2075 -593
rect 2041 -631 2075 -629
rect 2041 -703 2075 -697
rect 2041 -775 2075 -765
rect 2041 -847 2075 -833
rect 2041 -919 2075 -901
rect 2041 -991 2075 -969
rect 2041 -1063 2075 -1037
rect 2041 -1135 2075 -1105
rect 2041 -1207 2075 -1173
rect 2041 -1275 2075 -1241
rect 2041 -1343 2075 -1313
rect 2041 -1411 2075 -1385
rect 2041 -1479 2075 -1457
rect 2041 -1547 2075 -1529
rect 2041 -1615 2075 -1601
rect 2041 -1683 2075 -1673
rect 2041 -1751 2075 -1745
rect 2041 -1819 2075 -1817
rect 2041 -1855 2075 -1853
rect 2041 -1927 2075 -1921
rect 2041 -1999 2075 -1989
rect 2041 -2071 2075 -2057
rect 2041 -2143 2075 -2125
rect 2041 -2215 2075 -2193
rect 2041 -2287 2075 -2261
rect 2041 -2359 2075 -2329
rect 2041 -2431 2075 -2397
rect 2041 -2504 2075 -2465
rect 4099 2465 4133 2504
rect 4099 2397 4133 2431
rect 4099 2329 4133 2359
rect 4099 2261 4133 2287
rect 4099 2193 4133 2215
rect 4099 2125 4133 2143
rect 4099 2057 4133 2071
rect 4099 1989 4133 1999
rect 4099 1921 4133 1927
rect 4099 1853 4133 1855
rect 4099 1817 4133 1819
rect 4099 1745 4133 1751
rect 4099 1673 4133 1683
rect 4099 1601 4133 1615
rect 4099 1529 4133 1547
rect 4099 1457 4133 1479
rect 4099 1385 4133 1411
rect 4099 1313 4133 1343
rect 4099 1241 4133 1275
rect 4099 1173 4133 1207
rect 4099 1105 4133 1135
rect 4099 1037 4133 1063
rect 4099 969 4133 991
rect 4099 901 4133 919
rect 4099 833 4133 847
rect 4099 765 4133 775
rect 4099 697 4133 703
rect 4099 629 4133 631
rect 4099 593 4133 595
rect 4099 521 4133 527
rect 4099 449 4133 459
rect 4099 377 4133 391
rect 4099 305 4133 323
rect 4099 233 4133 255
rect 4099 161 4133 187
rect 4099 89 4133 119
rect 4099 17 4133 51
rect 4099 -51 4133 -17
rect 4099 -119 4133 -89
rect 4099 -187 4133 -161
rect 4099 -255 4133 -233
rect 4099 -323 4133 -305
rect 4099 -391 4133 -377
rect 4099 -459 4133 -449
rect 4099 -527 4133 -521
rect 4099 -595 4133 -593
rect 4099 -631 4133 -629
rect 4099 -703 4133 -697
rect 4099 -775 4133 -765
rect 4099 -847 4133 -833
rect 4099 -919 4133 -901
rect 4099 -991 4133 -969
rect 4099 -1063 4133 -1037
rect 4099 -1135 4133 -1105
rect 4099 -1207 4133 -1173
rect 4099 -1275 4133 -1241
rect 4099 -1343 4133 -1313
rect 4099 -1411 4133 -1385
rect 4099 -1479 4133 -1457
rect 4099 -1547 4133 -1529
rect 4099 -1615 4133 -1601
rect 4099 -1683 4133 -1673
rect 4099 -1751 4133 -1745
rect 4099 -1819 4133 -1817
rect 4099 -1855 4133 -1853
rect 4099 -1927 4133 -1921
rect 4099 -1999 4133 -1989
rect 4099 -2071 4133 -2057
rect 4099 -2143 4133 -2125
rect 4099 -2215 4133 -2193
rect 4099 -2287 4133 -2261
rect 4099 -2359 4133 -2329
rect 4099 -2431 4133 -2397
rect 4099 -2504 4133 -2465
rect 4213 2499 4247 2533
rect 4213 2431 4247 2465
rect 4213 2363 4247 2397
rect 4213 2295 4247 2329
rect 4213 2227 4247 2261
rect 4213 2159 4247 2193
rect 4213 2091 4247 2125
rect 4213 2023 4247 2057
rect 4213 1955 4247 1989
rect 4213 1887 4247 1921
rect 4213 1819 4247 1853
rect 4213 1751 4247 1785
rect 4213 1683 4247 1717
rect 4213 1615 4247 1649
rect 4213 1547 4247 1581
rect 4213 1479 4247 1513
rect 4213 1411 4247 1445
rect 4213 1343 4247 1377
rect 4213 1275 4247 1309
rect 4213 1207 4247 1241
rect 4213 1139 4247 1173
rect 4213 1071 4247 1105
rect 4213 1003 4247 1037
rect 4213 935 4247 969
rect 4213 867 4247 901
rect 4213 799 4247 833
rect 4213 731 4247 765
rect 4213 663 4247 697
rect 4213 595 4247 629
rect 4213 527 4247 561
rect 4213 459 4247 493
rect 4213 391 4247 425
rect 4213 323 4247 357
rect 4213 255 4247 289
rect 4213 187 4247 221
rect 4213 119 4247 153
rect 4213 51 4247 85
rect 4213 -17 4247 17
rect 4213 -85 4247 -51
rect 4213 -153 4247 -119
rect 4213 -221 4247 -187
rect 4213 -289 4247 -255
rect 4213 -357 4247 -323
rect 4213 -425 4247 -391
rect 4213 -493 4247 -459
rect 4213 -561 4247 -527
rect 4213 -629 4247 -595
rect 4213 -697 4247 -663
rect 4213 -765 4247 -731
rect 4213 -833 4247 -799
rect 4213 -901 4247 -867
rect 4213 -969 4247 -935
rect 4213 -1037 4247 -1003
rect 4213 -1105 4247 -1071
rect 4213 -1173 4247 -1139
rect 4213 -1241 4247 -1207
rect 4213 -1309 4247 -1275
rect 4213 -1377 4247 -1343
rect 4213 -1445 4247 -1411
rect 4213 -1513 4247 -1479
rect 4213 -1581 4247 -1547
rect 4213 -1649 4247 -1615
rect 4213 -1717 4247 -1683
rect 4213 -1785 4247 -1751
rect 4213 -1853 4247 -1819
rect 4213 -1921 4247 -1887
rect 4213 -1989 4247 -1955
rect 4213 -2057 4247 -2023
rect 4213 -2125 4247 -2091
rect 4213 -2193 4247 -2159
rect 4213 -2261 4247 -2227
rect 4213 -2329 4247 -2295
rect 4213 -2397 4247 -2363
rect 4213 -2465 4247 -2431
rect 4213 -2533 4247 -2499
rect -4247 -2640 -4213 -2567
rect -4087 -2572 -4056 -2538
rect -4006 -2572 -3988 -2538
rect -3934 -2572 -3920 -2538
rect -3862 -2572 -3852 -2538
rect -3790 -2572 -3784 -2538
rect -3718 -2572 -3716 -2538
rect -3682 -2572 -3680 -2538
rect -3614 -2572 -3608 -2538
rect -3546 -2572 -3536 -2538
rect -3478 -2572 -3464 -2538
rect -3410 -2572 -3392 -2538
rect -3342 -2572 -3320 -2538
rect -3274 -2572 -3248 -2538
rect -3206 -2572 -3176 -2538
rect -3138 -2572 -3104 -2538
rect -3070 -2572 -3036 -2538
rect -2998 -2572 -2968 -2538
rect -2926 -2572 -2900 -2538
rect -2854 -2572 -2832 -2538
rect -2782 -2572 -2764 -2538
rect -2710 -2572 -2696 -2538
rect -2638 -2572 -2628 -2538
rect -2566 -2572 -2560 -2538
rect -2494 -2572 -2492 -2538
rect -2458 -2572 -2456 -2538
rect -2390 -2572 -2384 -2538
rect -2322 -2572 -2312 -2538
rect -2254 -2572 -2240 -2538
rect -2186 -2572 -2168 -2538
rect -2118 -2572 -2087 -2538
rect -2029 -2572 -1998 -2538
rect -1948 -2572 -1930 -2538
rect -1876 -2572 -1862 -2538
rect -1804 -2572 -1794 -2538
rect -1732 -2572 -1726 -2538
rect -1660 -2572 -1658 -2538
rect -1624 -2572 -1622 -2538
rect -1556 -2572 -1550 -2538
rect -1488 -2572 -1478 -2538
rect -1420 -2572 -1406 -2538
rect -1352 -2572 -1334 -2538
rect -1284 -2572 -1262 -2538
rect -1216 -2572 -1190 -2538
rect -1148 -2572 -1118 -2538
rect -1080 -2572 -1046 -2538
rect -1012 -2572 -978 -2538
rect -940 -2572 -910 -2538
rect -868 -2572 -842 -2538
rect -796 -2572 -774 -2538
rect -724 -2572 -706 -2538
rect -652 -2572 -638 -2538
rect -580 -2572 -570 -2538
rect -508 -2572 -502 -2538
rect -436 -2572 -434 -2538
rect -400 -2572 -398 -2538
rect -332 -2572 -326 -2538
rect -264 -2572 -254 -2538
rect -196 -2572 -182 -2538
rect -128 -2572 -110 -2538
rect -60 -2572 -29 -2538
rect 29 -2572 60 -2538
rect 110 -2572 128 -2538
rect 182 -2572 196 -2538
rect 254 -2572 264 -2538
rect 326 -2572 332 -2538
rect 398 -2572 400 -2538
rect 434 -2572 436 -2538
rect 502 -2572 508 -2538
rect 570 -2572 580 -2538
rect 638 -2572 652 -2538
rect 706 -2572 724 -2538
rect 774 -2572 796 -2538
rect 842 -2572 868 -2538
rect 910 -2572 940 -2538
rect 978 -2572 1012 -2538
rect 1046 -2572 1080 -2538
rect 1118 -2572 1148 -2538
rect 1190 -2572 1216 -2538
rect 1262 -2572 1284 -2538
rect 1334 -2572 1352 -2538
rect 1406 -2572 1420 -2538
rect 1478 -2572 1488 -2538
rect 1550 -2572 1556 -2538
rect 1622 -2572 1624 -2538
rect 1658 -2572 1660 -2538
rect 1726 -2572 1732 -2538
rect 1794 -2572 1804 -2538
rect 1862 -2572 1876 -2538
rect 1930 -2572 1948 -2538
rect 1998 -2572 2029 -2538
rect 2087 -2572 2118 -2538
rect 2168 -2572 2186 -2538
rect 2240 -2572 2254 -2538
rect 2312 -2572 2322 -2538
rect 2384 -2572 2390 -2538
rect 2456 -2572 2458 -2538
rect 2492 -2572 2494 -2538
rect 2560 -2572 2566 -2538
rect 2628 -2572 2638 -2538
rect 2696 -2572 2710 -2538
rect 2764 -2572 2782 -2538
rect 2832 -2572 2854 -2538
rect 2900 -2572 2926 -2538
rect 2968 -2572 2998 -2538
rect 3036 -2572 3070 -2538
rect 3104 -2572 3138 -2538
rect 3176 -2572 3206 -2538
rect 3248 -2572 3274 -2538
rect 3320 -2572 3342 -2538
rect 3392 -2572 3410 -2538
rect 3464 -2572 3478 -2538
rect 3536 -2572 3546 -2538
rect 3608 -2572 3614 -2538
rect 3680 -2572 3682 -2538
rect 3716 -2572 3718 -2538
rect 3784 -2572 3790 -2538
rect 3852 -2572 3862 -2538
rect 3920 -2572 3934 -2538
rect 3988 -2572 4006 -2538
rect 4056 -2572 4087 -2538
rect 4213 -2640 4247 -2567
rect -4247 -2674 -4131 -2640
rect -4097 -2674 -4063 -2640
rect -4029 -2674 -3995 -2640
rect -3961 -2674 -3927 -2640
rect -3893 -2674 -3859 -2640
rect -3825 -2674 -3791 -2640
rect -3757 -2674 -3723 -2640
rect -3689 -2674 -3655 -2640
rect -3621 -2674 -3587 -2640
rect -3553 -2674 -3519 -2640
rect -3485 -2674 -3451 -2640
rect -3417 -2674 -3383 -2640
rect -3349 -2674 -3315 -2640
rect -3281 -2674 -3247 -2640
rect -3213 -2674 -3179 -2640
rect -3145 -2674 -3111 -2640
rect -3077 -2674 -3043 -2640
rect -3009 -2674 -2975 -2640
rect -2941 -2674 -2907 -2640
rect -2873 -2674 -2839 -2640
rect -2805 -2674 -2771 -2640
rect -2737 -2674 -2703 -2640
rect -2669 -2674 -2635 -2640
rect -2601 -2674 -2567 -2640
rect -2533 -2674 -2499 -2640
rect -2465 -2674 -2431 -2640
rect -2397 -2674 -2363 -2640
rect -2329 -2674 -2295 -2640
rect -2261 -2674 -2227 -2640
rect -2193 -2674 -2159 -2640
rect -2125 -2674 -2091 -2640
rect -2057 -2674 -2023 -2640
rect -1989 -2674 -1955 -2640
rect -1921 -2674 -1887 -2640
rect -1853 -2674 -1819 -2640
rect -1785 -2674 -1751 -2640
rect -1717 -2674 -1683 -2640
rect -1649 -2674 -1615 -2640
rect -1581 -2674 -1547 -2640
rect -1513 -2674 -1479 -2640
rect -1445 -2674 -1411 -2640
rect -1377 -2674 -1343 -2640
rect -1309 -2674 -1275 -2640
rect -1241 -2674 -1207 -2640
rect -1173 -2674 -1139 -2640
rect -1105 -2674 -1071 -2640
rect -1037 -2674 -1003 -2640
rect -969 -2674 -935 -2640
rect -901 -2674 -867 -2640
rect -833 -2674 -799 -2640
rect -765 -2674 -731 -2640
rect -697 -2674 -663 -2640
rect -629 -2674 -595 -2640
rect -561 -2674 -527 -2640
rect -493 -2674 -459 -2640
rect -425 -2674 -391 -2640
rect -357 -2674 -323 -2640
rect -289 -2674 -255 -2640
rect -221 -2674 -187 -2640
rect -153 -2674 -119 -2640
rect -85 -2674 -51 -2640
rect -17 -2674 17 -2640
rect 51 -2674 85 -2640
rect 119 -2674 153 -2640
rect 187 -2674 221 -2640
rect 255 -2674 289 -2640
rect 323 -2674 357 -2640
rect 391 -2674 425 -2640
rect 459 -2674 493 -2640
rect 527 -2674 561 -2640
rect 595 -2674 629 -2640
rect 663 -2674 697 -2640
rect 731 -2674 765 -2640
rect 799 -2674 833 -2640
rect 867 -2674 901 -2640
rect 935 -2674 969 -2640
rect 1003 -2674 1037 -2640
rect 1071 -2674 1105 -2640
rect 1139 -2674 1173 -2640
rect 1207 -2674 1241 -2640
rect 1275 -2674 1309 -2640
rect 1343 -2674 1377 -2640
rect 1411 -2674 1445 -2640
rect 1479 -2674 1513 -2640
rect 1547 -2674 1581 -2640
rect 1615 -2674 1649 -2640
rect 1683 -2674 1717 -2640
rect 1751 -2674 1785 -2640
rect 1819 -2674 1853 -2640
rect 1887 -2674 1921 -2640
rect 1955 -2674 1989 -2640
rect 2023 -2674 2057 -2640
rect 2091 -2674 2125 -2640
rect 2159 -2674 2193 -2640
rect 2227 -2674 2261 -2640
rect 2295 -2674 2329 -2640
rect 2363 -2674 2397 -2640
rect 2431 -2674 2465 -2640
rect 2499 -2674 2533 -2640
rect 2567 -2674 2601 -2640
rect 2635 -2674 2669 -2640
rect 2703 -2674 2737 -2640
rect 2771 -2674 2805 -2640
rect 2839 -2674 2873 -2640
rect 2907 -2674 2941 -2640
rect 2975 -2674 3009 -2640
rect 3043 -2674 3077 -2640
rect 3111 -2674 3145 -2640
rect 3179 -2674 3213 -2640
rect 3247 -2674 3281 -2640
rect 3315 -2674 3349 -2640
rect 3383 -2674 3417 -2640
rect 3451 -2674 3485 -2640
rect 3519 -2674 3553 -2640
rect 3587 -2674 3621 -2640
rect 3655 -2674 3689 -2640
rect 3723 -2674 3757 -2640
rect 3791 -2674 3825 -2640
rect 3859 -2674 3893 -2640
rect 3927 -2674 3961 -2640
rect 3995 -2674 4029 -2640
rect 4063 -2674 4097 -2640
rect 4131 -2674 4247 -2640
<< viali >>
rect -4040 2538 -4022 2572
rect -4022 2538 -4006 2572
rect -3968 2538 -3954 2572
rect -3954 2538 -3934 2572
rect -3896 2538 -3886 2572
rect -3886 2538 -3862 2572
rect -3824 2538 -3818 2572
rect -3818 2538 -3790 2572
rect -3752 2538 -3750 2572
rect -3750 2538 -3718 2572
rect -3680 2538 -3648 2572
rect -3648 2538 -3646 2572
rect -3608 2538 -3580 2572
rect -3580 2538 -3574 2572
rect -3536 2538 -3512 2572
rect -3512 2538 -3502 2572
rect -3464 2538 -3444 2572
rect -3444 2538 -3430 2572
rect -3392 2538 -3376 2572
rect -3376 2538 -3358 2572
rect -3320 2538 -3308 2572
rect -3308 2538 -3286 2572
rect -3248 2538 -3240 2572
rect -3240 2538 -3214 2572
rect -3176 2538 -3172 2572
rect -3172 2538 -3142 2572
rect -3104 2538 -3070 2572
rect -3032 2538 -3002 2572
rect -3002 2538 -2998 2572
rect -2960 2538 -2934 2572
rect -2934 2538 -2926 2572
rect -2888 2538 -2866 2572
rect -2866 2538 -2854 2572
rect -2816 2538 -2798 2572
rect -2798 2538 -2782 2572
rect -2744 2538 -2730 2572
rect -2730 2538 -2710 2572
rect -2672 2538 -2662 2572
rect -2662 2538 -2638 2572
rect -2600 2538 -2594 2572
rect -2594 2538 -2566 2572
rect -2528 2538 -2526 2572
rect -2526 2538 -2494 2572
rect -2456 2538 -2424 2572
rect -2424 2538 -2422 2572
rect -2384 2538 -2356 2572
rect -2356 2538 -2350 2572
rect -2312 2538 -2288 2572
rect -2288 2538 -2278 2572
rect -2240 2538 -2220 2572
rect -2220 2538 -2206 2572
rect -2168 2538 -2152 2572
rect -2152 2538 -2134 2572
rect -1982 2538 -1964 2572
rect -1964 2538 -1948 2572
rect -1910 2538 -1896 2572
rect -1896 2538 -1876 2572
rect -1838 2538 -1828 2572
rect -1828 2538 -1804 2572
rect -1766 2538 -1760 2572
rect -1760 2538 -1732 2572
rect -1694 2538 -1692 2572
rect -1692 2538 -1660 2572
rect -1622 2538 -1590 2572
rect -1590 2538 -1588 2572
rect -1550 2538 -1522 2572
rect -1522 2538 -1516 2572
rect -1478 2538 -1454 2572
rect -1454 2538 -1444 2572
rect -1406 2538 -1386 2572
rect -1386 2538 -1372 2572
rect -1334 2538 -1318 2572
rect -1318 2538 -1300 2572
rect -1262 2538 -1250 2572
rect -1250 2538 -1228 2572
rect -1190 2538 -1182 2572
rect -1182 2538 -1156 2572
rect -1118 2538 -1114 2572
rect -1114 2538 -1084 2572
rect -1046 2538 -1012 2572
rect -974 2538 -944 2572
rect -944 2538 -940 2572
rect -902 2538 -876 2572
rect -876 2538 -868 2572
rect -830 2538 -808 2572
rect -808 2538 -796 2572
rect -758 2538 -740 2572
rect -740 2538 -724 2572
rect -686 2538 -672 2572
rect -672 2538 -652 2572
rect -614 2538 -604 2572
rect -604 2538 -580 2572
rect -542 2538 -536 2572
rect -536 2538 -508 2572
rect -470 2538 -468 2572
rect -468 2538 -436 2572
rect -398 2538 -366 2572
rect -366 2538 -364 2572
rect -326 2538 -298 2572
rect -298 2538 -292 2572
rect -254 2538 -230 2572
rect -230 2538 -220 2572
rect -182 2538 -162 2572
rect -162 2538 -148 2572
rect -110 2538 -94 2572
rect -94 2538 -76 2572
rect 76 2538 94 2572
rect 94 2538 110 2572
rect 148 2538 162 2572
rect 162 2538 182 2572
rect 220 2538 230 2572
rect 230 2538 254 2572
rect 292 2538 298 2572
rect 298 2538 326 2572
rect 364 2538 366 2572
rect 366 2538 398 2572
rect 436 2538 468 2572
rect 468 2538 470 2572
rect 508 2538 536 2572
rect 536 2538 542 2572
rect 580 2538 604 2572
rect 604 2538 614 2572
rect 652 2538 672 2572
rect 672 2538 686 2572
rect 724 2538 740 2572
rect 740 2538 758 2572
rect 796 2538 808 2572
rect 808 2538 830 2572
rect 868 2538 876 2572
rect 876 2538 902 2572
rect 940 2538 944 2572
rect 944 2538 974 2572
rect 1012 2538 1046 2572
rect 1084 2538 1114 2572
rect 1114 2538 1118 2572
rect 1156 2538 1182 2572
rect 1182 2538 1190 2572
rect 1228 2538 1250 2572
rect 1250 2538 1262 2572
rect 1300 2538 1318 2572
rect 1318 2538 1334 2572
rect 1372 2538 1386 2572
rect 1386 2538 1406 2572
rect 1444 2538 1454 2572
rect 1454 2538 1478 2572
rect 1516 2538 1522 2572
rect 1522 2538 1550 2572
rect 1588 2538 1590 2572
rect 1590 2538 1622 2572
rect 1660 2538 1692 2572
rect 1692 2538 1694 2572
rect 1732 2538 1760 2572
rect 1760 2538 1766 2572
rect 1804 2538 1828 2572
rect 1828 2538 1838 2572
rect 1876 2538 1896 2572
rect 1896 2538 1910 2572
rect 1948 2538 1964 2572
rect 1964 2538 1982 2572
rect 2134 2538 2152 2572
rect 2152 2538 2168 2572
rect 2206 2538 2220 2572
rect 2220 2538 2240 2572
rect 2278 2538 2288 2572
rect 2288 2538 2312 2572
rect 2350 2538 2356 2572
rect 2356 2538 2384 2572
rect 2422 2538 2424 2572
rect 2424 2538 2456 2572
rect 2494 2538 2526 2572
rect 2526 2538 2528 2572
rect 2566 2538 2594 2572
rect 2594 2538 2600 2572
rect 2638 2538 2662 2572
rect 2662 2538 2672 2572
rect 2710 2538 2730 2572
rect 2730 2538 2744 2572
rect 2782 2538 2798 2572
rect 2798 2538 2816 2572
rect 2854 2538 2866 2572
rect 2866 2538 2888 2572
rect 2926 2538 2934 2572
rect 2934 2538 2960 2572
rect 2998 2538 3002 2572
rect 3002 2538 3032 2572
rect 3070 2538 3104 2572
rect 3142 2538 3172 2572
rect 3172 2538 3176 2572
rect 3214 2538 3240 2572
rect 3240 2538 3248 2572
rect 3286 2538 3308 2572
rect 3308 2538 3320 2572
rect 3358 2538 3376 2572
rect 3376 2538 3392 2572
rect 3430 2538 3444 2572
rect 3444 2538 3464 2572
rect 3502 2538 3512 2572
rect 3512 2538 3536 2572
rect 3574 2538 3580 2572
rect 3580 2538 3608 2572
rect 3646 2538 3648 2572
rect 3648 2538 3680 2572
rect 3718 2538 3750 2572
rect 3750 2538 3752 2572
rect 3790 2538 3818 2572
rect 3818 2538 3824 2572
rect 3862 2538 3886 2572
rect 3886 2538 3896 2572
rect 3934 2538 3954 2572
rect 3954 2538 3968 2572
rect 4006 2538 4022 2572
rect 4022 2538 4040 2572
rect -4133 2431 -4099 2465
rect -4133 2363 -4099 2393
rect -4133 2359 -4099 2363
rect -4133 2295 -4099 2321
rect -4133 2287 -4099 2295
rect -4133 2227 -4099 2249
rect -4133 2215 -4099 2227
rect -4133 2159 -4099 2177
rect -4133 2143 -4099 2159
rect -4133 2091 -4099 2105
rect -4133 2071 -4099 2091
rect -4133 2023 -4099 2033
rect -4133 1999 -4099 2023
rect -4133 1955 -4099 1961
rect -4133 1927 -4099 1955
rect -4133 1887 -4099 1889
rect -4133 1855 -4099 1887
rect -4133 1785 -4099 1817
rect -4133 1783 -4099 1785
rect -4133 1717 -4099 1745
rect -4133 1711 -4099 1717
rect -4133 1649 -4099 1673
rect -4133 1639 -4099 1649
rect -4133 1581 -4099 1601
rect -4133 1567 -4099 1581
rect -4133 1513 -4099 1529
rect -4133 1495 -4099 1513
rect -4133 1445 -4099 1457
rect -4133 1423 -4099 1445
rect -4133 1377 -4099 1385
rect -4133 1351 -4099 1377
rect -4133 1309 -4099 1313
rect -4133 1279 -4099 1309
rect -4133 1207 -4099 1241
rect -4133 1139 -4099 1169
rect -4133 1135 -4099 1139
rect -4133 1071 -4099 1097
rect -4133 1063 -4099 1071
rect -4133 1003 -4099 1025
rect -4133 991 -4099 1003
rect -4133 935 -4099 953
rect -4133 919 -4099 935
rect -4133 867 -4099 881
rect -4133 847 -4099 867
rect -4133 799 -4099 809
rect -4133 775 -4099 799
rect -4133 731 -4099 737
rect -4133 703 -4099 731
rect -4133 663 -4099 665
rect -4133 631 -4099 663
rect -4133 561 -4099 593
rect -4133 559 -4099 561
rect -4133 493 -4099 521
rect -4133 487 -4099 493
rect -4133 425 -4099 449
rect -4133 415 -4099 425
rect -4133 357 -4099 377
rect -4133 343 -4099 357
rect -4133 289 -4099 305
rect -4133 271 -4099 289
rect -4133 221 -4099 233
rect -4133 199 -4099 221
rect -4133 153 -4099 161
rect -4133 127 -4099 153
rect -4133 85 -4099 89
rect -4133 55 -4099 85
rect -4133 -17 -4099 17
rect -4133 -85 -4099 -55
rect -4133 -89 -4099 -85
rect -4133 -153 -4099 -127
rect -4133 -161 -4099 -153
rect -4133 -221 -4099 -199
rect -4133 -233 -4099 -221
rect -4133 -289 -4099 -271
rect -4133 -305 -4099 -289
rect -4133 -357 -4099 -343
rect -4133 -377 -4099 -357
rect -4133 -425 -4099 -415
rect -4133 -449 -4099 -425
rect -4133 -493 -4099 -487
rect -4133 -521 -4099 -493
rect -4133 -561 -4099 -559
rect -4133 -593 -4099 -561
rect -4133 -663 -4099 -631
rect -4133 -665 -4099 -663
rect -4133 -731 -4099 -703
rect -4133 -737 -4099 -731
rect -4133 -799 -4099 -775
rect -4133 -809 -4099 -799
rect -4133 -867 -4099 -847
rect -4133 -881 -4099 -867
rect -4133 -935 -4099 -919
rect -4133 -953 -4099 -935
rect -4133 -1003 -4099 -991
rect -4133 -1025 -4099 -1003
rect -4133 -1071 -4099 -1063
rect -4133 -1097 -4099 -1071
rect -4133 -1139 -4099 -1135
rect -4133 -1169 -4099 -1139
rect -4133 -1241 -4099 -1207
rect -4133 -1309 -4099 -1279
rect -4133 -1313 -4099 -1309
rect -4133 -1377 -4099 -1351
rect -4133 -1385 -4099 -1377
rect -4133 -1445 -4099 -1423
rect -4133 -1457 -4099 -1445
rect -4133 -1513 -4099 -1495
rect -4133 -1529 -4099 -1513
rect -4133 -1581 -4099 -1567
rect -4133 -1601 -4099 -1581
rect -4133 -1649 -4099 -1639
rect -4133 -1673 -4099 -1649
rect -4133 -1717 -4099 -1711
rect -4133 -1745 -4099 -1717
rect -4133 -1785 -4099 -1783
rect -4133 -1817 -4099 -1785
rect -4133 -1887 -4099 -1855
rect -4133 -1889 -4099 -1887
rect -4133 -1955 -4099 -1927
rect -4133 -1961 -4099 -1955
rect -4133 -2023 -4099 -1999
rect -4133 -2033 -4099 -2023
rect -4133 -2091 -4099 -2071
rect -4133 -2105 -4099 -2091
rect -4133 -2159 -4099 -2143
rect -4133 -2177 -4099 -2159
rect -4133 -2227 -4099 -2215
rect -4133 -2249 -4099 -2227
rect -4133 -2295 -4099 -2287
rect -4133 -2321 -4099 -2295
rect -4133 -2363 -4099 -2359
rect -4133 -2393 -4099 -2363
rect -4133 -2465 -4099 -2431
rect -2075 2431 -2041 2465
rect -2075 2363 -2041 2393
rect -2075 2359 -2041 2363
rect -2075 2295 -2041 2321
rect -2075 2287 -2041 2295
rect -2075 2227 -2041 2249
rect -2075 2215 -2041 2227
rect -2075 2159 -2041 2177
rect -2075 2143 -2041 2159
rect -2075 2091 -2041 2105
rect -2075 2071 -2041 2091
rect -2075 2023 -2041 2033
rect -2075 1999 -2041 2023
rect -2075 1955 -2041 1961
rect -2075 1927 -2041 1955
rect -2075 1887 -2041 1889
rect -2075 1855 -2041 1887
rect -2075 1785 -2041 1817
rect -2075 1783 -2041 1785
rect -2075 1717 -2041 1745
rect -2075 1711 -2041 1717
rect -2075 1649 -2041 1673
rect -2075 1639 -2041 1649
rect -2075 1581 -2041 1601
rect -2075 1567 -2041 1581
rect -2075 1513 -2041 1529
rect -2075 1495 -2041 1513
rect -2075 1445 -2041 1457
rect -2075 1423 -2041 1445
rect -2075 1377 -2041 1385
rect -2075 1351 -2041 1377
rect -2075 1309 -2041 1313
rect -2075 1279 -2041 1309
rect -2075 1207 -2041 1241
rect -2075 1139 -2041 1169
rect -2075 1135 -2041 1139
rect -2075 1071 -2041 1097
rect -2075 1063 -2041 1071
rect -2075 1003 -2041 1025
rect -2075 991 -2041 1003
rect -2075 935 -2041 953
rect -2075 919 -2041 935
rect -2075 867 -2041 881
rect -2075 847 -2041 867
rect -2075 799 -2041 809
rect -2075 775 -2041 799
rect -2075 731 -2041 737
rect -2075 703 -2041 731
rect -2075 663 -2041 665
rect -2075 631 -2041 663
rect -2075 561 -2041 593
rect -2075 559 -2041 561
rect -2075 493 -2041 521
rect -2075 487 -2041 493
rect -2075 425 -2041 449
rect -2075 415 -2041 425
rect -2075 357 -2041 377
rect -2075 343 -2041 357
rect -2075 289 -2041 305
rect -2075 271 -2041 289
rect -2075 221 -2041 233
rect -2075 199 -2041 221
rect -2075 153 -2041 161
rect -2075 127 -2041 153
rect -2075 85 -2041 89
rect -2075 55 -2041 85
rect -2075 -17 -2041 17
rect -2075 -85 -2041 -55
rect -2075 -89 -2041 -85
rect -2075 -153 -2041 -127
rect -2075 -161 -2041 -153
rect -2075 -221 -2041 -199
rect -2075 -233 -2041 -221
rect -2075 -289 -2041 -271
rect -2075 -305 -2041 -289
rect -2075 -357 -2041 -343
rect -2075 -377 -2041 -357
rect -2075 -425 -2041 -415
rect -2075 -449 -2041 -425
rect -2075 -493 -2041 -487
rect -2075 -521 -2041 -493
rect -2075 -561 -2041 -559
rect -2075 -593 -2041 -561
rect -2075 -663 -2041 -631
rect -2075 -665 -2041 -663
rect -2075 -731 -2041 -703
rect -2075 -737 -2041 -731
rect -2075 -799 -2041 -775
rect -2075 -809 -2041 -799
rect -2075 -867 -2041 -847
rect -2075 -881 -2041 -867
rect -2075 -935 -2041 -919
rect -2075 -953 -2041 -935
rect -2075 -1003 -2041 -991
rect -2075 -1025 -2041 -1003
rect -2075 -1071 -2041 -1063
rect -2075 -1097 -2041 -1071
rect -2075 -1139 -2041 -1135
rect -2075 -1169 -2041 -1139
rect -2075 -1241 -2041 -1207
rect -2075 -1309 -2041 -1279
rect -2075 -1313 -2041 -1309
rect -2075 -1377 -2041 -1351
rect -2075 -1385 -2041 -1377
rect -2075 -1445 -2041 -1423
rect -2075 -1457 -2041 -1445
rect -2075 -1513 -2041 -1495
rect -2075 -1529 -2041 -1513
rect -2075 -1581 -2041 -1567
rect -2075 -1601 -2041 -1581
rect -2075 -1649 -2041 -1639
rect -2075 -1673 -2041 -1649
rect -2075 -1717 -2041 -1711
rect -2075 -1745 -2041 -1717
rect -2075 -1785 -2041 -1783
rect -2075 -1817 -2041 -1785
rect -2075 -1887 -2041 -1855
rect -2075 -1889 -2041 -1887
rect -2075 -1955 -2041 -1927
rect -2075 -1961 -2041 -1955
rect -2075 -2023 -2041 -1999
rect -2075 -2033 -2041 -2023
rect -2075 -2091 -2041 -2071
rect -2075 -2105 -2041 -2091
rect -2075 -2159 -2041 -2143
rect -2075 -2177 -2041 -2159
rect -2075 -2227 -2041 -2215
rect -2075 -2249 -2041 -2227
rect -2075 -2295 -2041 -2287
rect -2075 -2321 -2041 -2295
rect -2075 -2363 -2041 -2359
rect -2075 -2393 -2041 -2363
rect -2075 -2465 -2041 -2431
rect -17 2431 17 2465
rect -17 2363 17 2393
rect -17 2359 17 2363
rect -17 2295 17 2321
rect -17 2287 17 2295
rect -17 2227 17 2249
rect -17 2215 17 2227
rect -17 2159 17 2177
rect -17 2143 17 2159
rect -17 2091 17 2105
rect -17 2071 17 2091
rect -17 2023 17 2033
rect -17 1999 17 2023
rect -17 1955 17 1961
rect -17 1927 17 1955
rect -17 1887 17 1889
rect -17 1855 17 1887
rect -17 1785 17 1817
rect -17 1783 17 1785
rect -17 1717 17 1745
rect -17 1711 17 1717
rect -17 1649 17 1673
rect -17 1639 17 1649
rect -17 1581 17 1601
rect -17 1567 17 1581
rect -17 1513 17 1529
rect -17 1495 17 1513
rect -17 1445 17 1457
rect -17 1423 17 1445
rect -17 1377 17 1385
rect -17 1351 17 1377
rect -17 1309 17 1313
rect -17 1279 17 1309
rect -17 1207 17 1241
rect -17 1139 17 1169
rect -17 1135 17 1139
rect -17 1071 17 1097
rect -17 1063 17 1071
rect -17 1003 17 1025
rect -17 991 17 1003
rect -17 935 17 953
rect -17 919 17 935
rect -17 867 17 881
rect -17 847 17 867
rect -17 799 17 809
rect -17 775 17 799
rect -17 731 17 737
rect -17 703 17 731
rect -17 663 17 665
rect -17 631 17 663
rect -17 561 17 593
rect -17 559 17 561
rect -17 493 17 521
rect -17 487 17 493
rect -17 425 17 449
rect -17 415 17 425
rect -17 357 17 377
rect -17 343 17 357
rect -17 289 17 305
rect -17 271 17 289
rect -17 221 17 233
rect -17 199 17 221
rect -17 153 17 161
rect -17 127 17 153
rect -17 85 17 89
rect -17 55 17 85
rect -17 -17 17 17
rect -17 -85 17 -55
rect -17 -89 17 -85
rect -17 -153 17 -127
rect -17 -161 17 -153
rect -17 -221 17 -199
rect -17 -233 17 -221
rect -17 -289 17 -271
rect -17 -305 17 -289
rect -17 -357 17 -343
rect -17 -377 17 -357
rect -17 -425 17 -415
rect -17 -449 17 -425
rect -17 -493 17 -487
rect -17 -521 17 -493
rect -17 -561 17 -559
rect -17 -593 17 -561
rect -17 -663 17 -631
rect -17 -665 17 -663
rect -17 -731 17 -703
rect -17 -737 17 -731
rect -17 -799 17 -775
rect -17 -809 17 -799
rect -17 -867 17 -847
rect -17 -881 17 -867
rect -17 -935 17 -919
rect -17 -953 17 -935
rect -17 -1003 17 -991
rect -17 -1025 17 -1003
rect -17 -1071 17 -1063
rect -17 -1097 17 -1071
rect -17 -1139 17 -1135
rect -17 -1169 17 -1139
rect -17 -1241 17 -1207
rect -17 -1309 17 -1279
rect -17 -1313 17 -1309
rect -17 -1377 17 -1351
rect -17 -1385 17 -1377
rect -17 -1445 17 -1423
rect -17 -1457 17 -1445
rect -17 -1513 17 -1495
rect -17 -1529 17 -1513
rect -17 -1581 17 -1567
rect -17 -1601 17 -1581
rect -17 -1649 17 -1639
rect -17 -1673 17 -1649
rect -17 -1717 17 -1711
rect -17 -1745 17 -1717
rect -17 -1785 17 -1783
rect -17 -1817 17 -1785
rect -17 -1887 17 -1855
rect -17 -1889 17 -1887
rect -17 -1955 17 -1927
rect -17 -1961 17 -1955
rect -17 -2023 17 -1999
rect -17 -2033 17 -2023
rect -17 -2091 17 -2071
rect -17 -2105 17 -2091
rect -17 -2159 17 -2143
rect -17 -2177 17 -2159
rect -17 -2227 17 -2215
rect -17 -2249 17 -2227
rect -17 -2295 17 -2287
rect -17 -2321 17 -2295
rect -17 -2363 17 -2359
rect -17 -2393 17 -2363
rect -17 -2465 17 -2431
rect 2041 2431 2075 2465
rect 2041 2363 2075 2393
rect 2041 2359 2075 2363
rect 2041 2295 2075 2321
rect 2041 2287 2075 2295
rect 2041 2227 2075 2249
rect 2041 2215 2075 2227
rect 2041 2159 2075 2177
rect 2041 2143 2075 2159
rect 2041 2091 2075 2105
rect 2041 2071 2075 2091
rect 2041 2023 2075 2033
rect 2041 1999 2075 2023
rect 2041 1955 2075 1961
rect 2041 1927 2075 1955
rect 2041 1887 2075 1889
rect 2041 1855 2075 1887
rect 2041 1785 2075 1817
rect 2041 1783 2075 1785
rect 2041 1717 2075 1745
rect 2041 1711 2075 1717
rect 2041 1649 2075 1673
rect 2041 1639 2075 1649
rect 2041 1581 2075 1601
rect 2041 1567 2075 1581
rect 2041 1513 2075 1529
rect 2041 1495 2075 1513
rect 2041 1445 2075 1457
rect 2041 1423 2075 1445
rect 2041 1377 2075 1385
rect 2041 1351 2075 1377
rect 2041 1309 2075 1313
rect 2041 1279 2075 1309
rect 2041 1207 2075 1241
rect 2041 1139 2075 1169
rect 2041 1135 2075 1139
rect 2041 1071 2075 1097
rect 2041 1063 2075 1071
rect 2041 1003 2075 1025
rect 2041 991 2075 1003
rect 2041 935 2075 953
rect 2041 919 2075 935
rect 2041 867 2075 881
rect 2041 847 2075 867
rect 2041 799 2075 809
rect 2041 775 2075 799
rect 2041 731 2075 737
rect 2041 703 2075 731
rect 2041 663 2075 665
rect 2041 631 2075 663
rect 2041 561 2075 593
rect 2041 559 2075 561
rect 2041 493 2075 521
rect 2041 487 2075 493
rect 2041 425 2075 449
rect 2041 415 2075 425
rect 2041 357 2075 377
rect 2041 343 2075 357
rect 2041 289 2075 305
rect 2041 271 2075 289
rect 2041 221 2075 233
rect 2041 199 2075 221
rect 2041 153 2075 161
rect 2041 127 2075 153
rect 2041 85 2075 89
rect 2041 55 2075 85
rect 2041 -17 2075 17
rect 2041 -85 2075 -55
rect 2041 -89 2075 -85
rect 2041 -153 2075 -127
rect 2041 -161 2075 -153
rect 2041 -221 2075 -199
rect 2041 -233 2075 -221
rect 2041 -289 2075 -271
rect 2041 -305 2075 -289
rect 2041 -357 2075 -343
rect 2041 -377 2075 -357
rect 2041 -425 2075 -415
rect 2041 -449 2075 -425
rect 2041 -493 2075 -487
rect 2041 -521 2075 -493
rect 2041 -561 2075 -559
rect 2041 -593 2075 -561
rect 2041 -663 2075 -631
rect 2041 -665 2075 -663
rect 2041 -731 2075 -703
rect 2041 -737 2075 -731
rect 2041 -799 2075 -775
rect 2041 -809 2075 -799
rect 2041 -867 2075 -847
rect 2041 -881 2075 -867
rect 2041 -935 2075 -919
rect 2041 -953 2075 -935
rect 2041 -1003 2075 -991
rect 2041 -1025 2075 -1003
rect 2041 -1071 2075 -1063
rect 2041 -1097 2075 -1071
rect 2041 -1139 2075 -1135
rect 2041 -1169 2075 -1139
rect 2041 -1241 2075 -1207
rect 2041 -1309 2075 -1279
rect 2041 -1313 2075 -1309
rect 2041 -1377 2075 -1351
rect 2041 -1385 2075 -1377
rect 2041 -1445 2075 -1423
rect 2041 -1457 2075 -1445
rect 2041 -1513 2075 -1495
rect 2041 -1529 2075 -1513
rect 2041 -1581 2075 -1567
rect 2041 -1601 2075 -1581
rect 2041 -1649 2075 -1639
rect 2041 -1673 2075 -1649
rect 2041 -1717 2075 -1711
rect 2041 -1745 2075 -1717
rect 2041 -1785 2075 -1783
rect 2041 -1817 2075 -1785
rect 2041 -1887 2075 -1855
rect 2041 -1889 2075 -1887
rect 2041 -1955 2075 -1927
rect 2041 -1961 2075 -1955
rect 2041 -2023 2075 -1999
rect 2041 -2033 2075 -2023
rect 2041 -2091 2075 -2071
rect 2041 -2105 2075 -2091
rect 2041 -2159 2075 -2143
rect 2041 -2177 2075 -2159
rect 2041 -2227 2075 -2215
rect 2041 -2249 2075 -2227
rect 2041 -2295 2075 -2287
rect 2041 -2321 2075 -2295
rect 2041 -2363 2075 -2359
rect 2041 -2393 2075 -2363
rect 2041 -2465 2075 -2431
rect 4099 2431 4133 2465
rect 4099 2363 4133 2393
rect 4099 2359 4133 2363
rect 4099 2295 4133 2321
rect 4099 2287 4133 2295
rect 4099 2227 4133 2249
rect 4099 2215 4133 2227
rect 4099 2159 4133 2177
rect 4099 2143 4133 2159
rect 4099 2091 4133 2105
rect 4099 2071 4133 2091
rect 4099 2023 4133 2033
rect 4099 1999 4133 2023
rect 4099 1955 4133 1961
rect 4099 1927 4133 1955
rect 4099 1887 4133 1889
rect 4099 1855 4133 1887
rect 4099 1785 4133 1817
rect 4099 1783 4133 1785
rect 4099 1717 4133 1745
rect 4099 1711 4133 1717
rect 4099 1649 4133 1673
rect 4099 1639 4133 1649
rect 4099 1581 4133 1601
rect 4099 1567 4133 1581
rect 4099 1513 4133 1529
rect 4099 1495 4133 1513
rect 4099 1445 4133 1457
rect 4099 1423 4133 1445
rect 4099 1377 4133 1385
rect 4099 1351 4133 1377
rect 4099 1309 4133 1313
rect 4099 1279 4133 1309
rect 4099 1207 4133 1241
rect 4099 1139 4133 1169
rect 4099 1135 4133 1139
rect 4099 1071 4133 1097
rect 4099 1063 4133 1071
rect 4099 1003 4133 1025
rect 4099 991 4133 1003
rect 4099 935 4133 953
rect 4099 919 4133 935
rect 4099 867 4133 881
rect 4099 847 4133 867
rect 4099 799 4133 809
rect 4099 775 4133 799
rect 4099 731 4133 737
rect 4099 703 4133 731
rect 4099 663 4133 665
rect 4099 631 4133 663
rect 4099 561 4133 593
rect 4099 559 4133 561
rect 4099 493 4133 521
rect 4099 487 4133 493
rect 4099 425 4133 449
rect 4099 415 4133 425
rect 4099 357 4133 377
rect 4099 343 4133 357
rect 4099 289 4133 305
rect 4099 271 4133 289
rect 4099 221 4133 233
rect 4099 199 4133 221
rect 4099 153 4133 161
rect 4099 127 4133 153
rect 4099 85 4133 89
rect 4099 55 4133 85
rect 4099 -17 4133 17
rect 4099 -85 4133 -55
rect 4099 -89 4133 -85
rect 4099 -153 4133 -127
rect 4099 -161 4133 -153
rect 4099 -221 4133 -199
rect 4099 -233 4133 -221
rect 4099 -289 4133 -271
rect 4099 -305 4133 -289
rect 4099 -357 4133 -343
rect 4099 -377 4133 -357
rect 4099 -425 4133 -415
rect 4099 -449 4133 -425
rect 4099 -493 4133 -487
rect 4099 -521 4133 -493
rect 4099 -561 4133 -559
rect 4099 -593 4133 -561
rect 4099 -663 4133 -631
rect 4099 -665 4133 -663
rect 4099 -731 4133 -703
rect 4099 -737 4133 -731
rect 4099 -799 4133 -775
rect 4099 -809 4133 -799
rect 4099 -867 4133 -847
rect 4099 -881 4133 -867
rect 4099 -935 4133 -919
rect 4099 -953 4133 -935
rect 4099 -1003 4133 -991
rect 4099 -1025 4133 -1003
rect 4099 -1071 4133 -1063
rect 4099 -1097 4133 -1071
rect 4099 -1139 4133 -1135
rect 4099 -1169 4133 -1139
rect 4099 -1241 4133 -1207
rect 4099 -1309 4133 -1279
rect 4099 -1313 4133 -1309
rect 4099 -1377 4133 -1351
rect 4099 -1385 4133 -1377
rect 4099 -1445 4133 -1423
rect 4099 -1457 4133 -1445
rect 4099 -1513 4133 -1495
rect 4099 -1529 4133 -1513
rect 4099 -1581 4133 -1567
rect 4099 -1601 4133 -1581
rect 4099 -1649 4133 -1639
rect 4099 -1673 4133 -1649
rect 4099 -1717 4133 -1711
rect 4099 -1745 4133 -1717
rect 4099 -1785 4133 -1783
rect 4099 -1817 4133 -1785
rect 4099 -1887 4133 -1855
rect 4099 -1889 4133 -1887
rect 4099 -1955 4133 -1927
rect 4099 -1961 4133 -1955
rect 4099 -2023 4133 -1999
rect 4099 -2033 4133 -2023
rect 4099 -2091 4133 -2071
rect 4099 -2105 4133 -2091
rect 4099 -2159 4133 -2143
rect 4099 -2177 4133 -2159
rect 4099 -2227 4133 -2215
rect 4099 -2249 4133 -2227
rect 4099 -2295 4133 -2287
rect 4099 -2321 4133 -2295
rect 4099 -2363 4133 -2359
rect 4099 -2393 4133 -2363
rect 4099 -2465 4133 -2431
rect -4040 -2572 -4022 -2538
rect -4022 -2572 -4006 -2538
rect -3968 -2572 -3954 -2538
rect -3954 -2572 -3934 -2538
rect -3896 -2572 -3886 -2538
rect -3886 -2572 -3862 -2538
rect -3824 -2572 -3818 -2538
rect -3818 -2572 -3790 -2538
rect -3752 -2572 -3750 -2538
rect -3750 -2572 -3718 -2538
rect -3680 -2572 -3648 -2538
rect -3648 -2572 -3646 -2538
rect -3608 -2572 -3580 -2538
rect -3580 -2572 -3574 -2538
rect -3536 -2572 -3512 -2538
rect -3512 -2572 -3502 -2538
rect -3464 -2572 -3444 -2538
rect -3444 -2572 -3430 -2538
rect -3392 -2572 -3376 -2538
rect -3376 -2572 -3358 -2538
rect -3320 -2572 -3308 -2538
rect -3308 -2572 -3286 -2538
rect -3248 -2572 -3240 -2538
rect -3240 -2572 -3214 -2538
rect -3176 -2572 -3172 -2538
rect -3172 -2572 -3142 -2538
rect -3104 -2572 -3070 -2538
rect -3032 -2572 -3002 -2538
rect -3002 -2572 -2998 -2538
rect -2960 -2572 -2934 -2538
rect -2934 -2572 -2926 -2538
rect -2888 -2572 -2866 -2538
rect -2866 -2572 -2854 -2538
rect -2816 -2572 -2798 -2538
rect -2798 -2572 -2782 -2538
rect -2744 -2572 -2730 -2538
rect -2730 -2572 -2710 -2538
rect -2672 -2572 -2662 -2538
rect -2662 -2572 -2638 -2538
rect -2600 -2572 -2594 -2538
rect -2594 -2572 -2566 -2538
rect -2528 -2572 -2526 -2538
rect -2526 -2572 -2494 -2538
rect -2456 -2572 -2424 -2538
rect -2424 -2572 -2422 -2538
rect -2384 -2572 -2356 -2538
rect -2356 -2572 -2350 -2538
rect -2312 -2572 -2288 -2538
rect -2288 -2572 -2278 -2538
rect -2240 -2572 -2220 -2538
rect -2220 -2572 -2206 -2538
rect -2168 -2572 -2152 -2538
rect -2152 -2572 -2134 -2538
rect -1982 -2572 -1964 -2538
rect -1964 -2572 -1948 -2538
rect -1910 -2572 -1896 -2538
rect -1896 -2572 -1876 -2538
rect -1838 -2572 -1828 -2538
rect -1828 -2572 -1804 -2538
rect -1766 -2572 -1760 -2538
rect -1760 -2572 -1732 -2538
rect -1694 -2572 -1692 -2538
rect -1692 -2572 -1660 -2538
rect -1622 -2572 -1590 -2538
rect -1590 -2572 -1588 -2538
rect -1550 -2572 -1522 -2538
rect -1522 -2572 -1516 -2538
rect -1478 -2572 -1454 -2538
rect -1454 -2572 -1444 -2538
rect -1406 -2572 -1386 -2538
rect -1386 -2572 -1372 -2538
rect -1334 -2572 -1318 -2538
rect -1318 -2572 -1300 -2538
rect -1262 -2572 -1250 -2538
rect -1250 -2572 -1228 -2538
rect -1190 -2572 -1182 -2538
rect -1182 -2572 -1156 -2538
rect -1118 -2572 -1114 -2538
rect -1114 -2572 -1084 -2538
rect -1046 -2572 -1012 -2538
rect -974 -2572 -944 -2538
rect -944 -2572 -940 -2538
rect -902 -2572 -876 -2538
rect -876 -2572 -868 -2538
rect -830 -2572 -808 -2538
rect -808 -2572 -796 -2538
rect -758 -2572 -740 -2538
rect -740 -2572 -724 -2538
rect -686 -2572 -672 -2538
rect -672 -2572 -652 -2538
rect -614 -2572 -604 -2538
rect -604 -2572 -580 -2538
rect -542 -2572 -536 -2538
rect -536 -2572 -508 -2538
rect -470 -2572 -468 -2538
rect -468 -2572 -436 -2538
rect -398 -2572 -366 -2538
rect -366 -2572 -364 -2538
rect -326 -2572 -298 -2538
rect -298 -2572 -292 -2538
rect -254 -2572 -230 -2538
rect -230 -2572 -220 -2538
rect -182 -2572 -162 -2538
rect -162 -2572 -148 -2538
rect -110 -2572 -94 -2538
rect -94 -2572 -76 -2538
rect 76 -2572 94 -2538
rect 94 -2572 110 -2538
rect 148 -2572 162 -2538
rect 162 -2572 182 -2538
rect 220 -2572 230 -2538
rect 230 -2572 254 -2538
rect 292 -2572 298 -2538
rect 298 -2572 326 -2538
rect 364 -2572 366 -2538
rect 366 -2572 398 -2538
rect 436 -2572 468 -2538
rect 468 -2572 470 -2538
rect 508 -2572 536 -2538
rect 536 -2572 542 -2538
rect 580 -2572 604 -2538
rect 604 -2572 614 -2538
rect 652 -2572 672 -2538
rect 672 -2572 686 -2538
rect 724 -2572 740 -2538
rect 740 -2572 758 -2538
rect 796 -2572 808 -2538
rect 808 -2572 830 -2538
rect 868 -2572 876 -2538
rect 876 -2572 902 -2538
rect 940 -2572 944 -2538
rect 944 -2572 974 -2538
rect 1012 -2572 1046 -2538
rect 1084 -2572 1114 -2538
rect 1114 -2572 1118 -2538
rect 1156 -2572 1182 -2538
rect 1182 -2572 1190 -2538
rect 1228 -2572 1250 -2538
rect 1250 -2572 1262 -2538
rect 1300 -2572 1318 -2538
rect 1318 -2572 1334 -2538
rect 1372 -2572 1386 -2538
rect 1386 -2572 1406 -2538
rect 1444 -2572 1454 -2538
rect 1454 -2572 1478 -2538
rect 1516 -2572 1522 -2538
rect 1522 -2572 1550 -2538
rect 1588 -2572 1590 -2538
rect 1590 -2572 1622 -2538
rect 1660 -2572 1692 -2538
rect 1692 -2572 1694 -2538
rect 1732 -2572 1760 -2538
rect 1760 -2572 1766 -2538
rect 1804 -2572 1828 -2538
rect 1828 -2572 1838 -2538
rect 1876 -2572 1896 -2538
rect 1896 -2572 1910 -2538
rect 1948 -2572 1964 -2538
rect 1964 -2572 1982 -2538
rect 2134 -2572 2152 -2538
rect 2152 -2572 2168 -2538
rect 2206 -2572 2220 -2538
rect 2220 -2572 2240 -2538
rect 2278 -2572 2288 -2538
rect 2288 -2572 2312 -2538
rect 2350 -2572 2356 -2538
rect 2356 -2572 2384 -2538
rect 2422 -2572 2424 -2538
rect 2424 -2572 2456 -2538
rect 2494 -2572 2526 -2538
rect 2526 -2572 2528 -2538
rect 2566 -2572 2594 -2538
rect 2594 -2572 2600 -2538
rect 2638 -2572 2662 -2538
rect 2662 -2572 2672 -2538
rect 2710 -2572 2730 -2538
rect 2730 -2572 2744 -2538
rect 2782 -2572 2798 -2538
rect 2798 -2572 2816 -2538
rect 2854 -2572 2866 -2538
rect 2866 -2572 2888 -2538
rect 2926 -2572 2934 -2538
rect 2934 -2572 2960 -2538
rect 2998 -2572 3002 -2538
rect 3002 -2572 3032 -2538
rect 3070 -2572 3104 -2538
rect 3142 -2572 3172 -2538
rect 3172 -2572 3176 -2538
rect 3214 -2572 3240 -2538
rect 3240 -2572 3248 -2538
rect 3286 -2572 3308 -2538
rect 3308 -2572 3320 -2538
rect 3358 -2572 3376 -2538
rect 3376 -2572 3392 -2538
rect 3430 -2572 3444 -2538
rect 3444 -2572 3464 -2538
rect 3502 -2572 3512 -2538
rect 3512 -2572 3536 -2538
rect 3574 -2572 3580 -2538
rect 3580 -2572 3608 -2538
rect 3646 -2572 3648 -2538
rect 3648 -2572 3680 -2538
rect 3718 -2572 3750 -2538
rect 3750 -2572 3752 -2538
rect 3790 -2572 3818 -2538
rect 3818 -2572 3824 -2538
rect 3862 -2572 3886 -2538
rect 3886 -2572 3896 -2538
rect 3934 -2572 3954 -2538
rect 3954 -2572 3968 -2538
rect 4006 -2572 4022 -2538
rect 4022 -2572 4040 -2538
<< metal1 >>
rect -4083 2572 -2091 2578
rect -4083 2538 -4040 2572
rect -4006 2538 -3968 2572
rect -3934 2538 -3896 2572
rect -3862 2538 -3824 2572
rect -3790 2538 -3752 2572
rect -3718 2538 -3680 2572
rect -3646 2538 -3608 2572
rect -3574 2538 -3536 2572
rect -3502 2538 -3464 2572
rect -3430 2538 -3392 2572
rect -3358 2538 -3320 2572
rect -3286 2538 -3248 2572
rect -3214 2538 -3176 2572
rect -3142 2538 -3104 2572
rect -3070 2538 -3032 2572
rect -2998 2538 -2960 2572
rect -2926 2538 -2888 2572
rect -2854 2538 -2816 2572
rect -2782 2538 -2744 2572
rect -2710 2538 -2672 2572
rect -2638 2538 -2600 2572
rect -2566 2538 -2528 2572
rect -2494 2538 -2456 2572
rect -2422 2538 -2384 2572
rect -2350 2538 -2312 2572
rect -2278 2538 -2240 2572
rect -2206 2538 -2168 2572
rect -2134 2538 -2091 2572
rect -4083 2532 -2091 2538
rect -2025 2572 -33 2578
rect -2025 2538 -1982 2572
rect -1948 2538 -1910 2572
rect -1876 2538 -1838 2572
rect -1804 2538 -1766 2572
rect -1732 2538 -1694 2572
rect -1660 2538 -1622 2572
rect -1588 2538 -1550 2572
rect -1516 2538 -1478 2572
rect -1444 2538 -1406 2572
rect -1372 2538 -1334 2572
rect -1300 2538 -1262 2572
rect -1228 2538 -1190 2572
rect -1156 2538 -1118 2572
rect -1084 2538 -1046 2572
rect -1012 2538 -974 2572
rect -940 2538 -902 2572
rect -868 2538 -830 2572
rect -796 2538 -758 2572
rect -724 2538 -686 2572
rect -652 2538 -614 2572
rect -580 2538 -542 2572
rect -508 2538 -470 2572
rect -436 2538 -398 2572
rect -364 2538 -326 2572
rect -292 2538 -254 2572
rect -220 2538 -182 2572
rect -148 2538 -110 2572
rect -76 2538 -33 2572
rect -2025 2532 -33 2538
rect 33 2572 2025 2578
rect 33 2538 76 2572
rect 110 2538 148 2572
rect 182 2538 220 2572
rect 254 2538 292 2572
rect 326 2538 364 2572
rect 398 2538 436 2572
rect 470 2538 508 2572
rect 542 2538 580 2572
rect 614 2538 652 2572
rect 686 2538 724 2572
rect 758 2538 796 2572
rect 830 2538 868 2572
rect 902 2538 940 2572
rect 974 2538 1012 2572
rect 1046 2538 1084 2572
rect 1118 2538 1156 2572
rect 1190 2538 1228 2572
rect 1262 2538 1300 2572
rect 1334 2538 1372 2572
rect 1406 2538 1444 2572
rect 1478 2538 1516 2572
rect 1550 2538 1588 2572
rect 1622 2538 1660 2572
rect 1694 2538 1732 2572
rect 1766 2538 1804 2572
rect 1838 2538 1876 2572
rect 1910 2538 1948 2572
rect 1982 2538 2025 2572
rect 33 2532 2025 2538
rect 2091 2572 4083 2578
rect 2091 2538 2134 2572
rect 2168 2538 2206 2572
rect 2240 2538 2278 2572
rect 2312 2538 2350 2572
rect 2384 2538 2422 2572
rect 2456 2538 2494 2572
rect 2528 2538 2566 2572
rect 2600 2538 2638 2572
rect 2672 2538 2710 2572
rect 2744 2538 2782 2572
rect 2816 2538 2854 2572
rect 2888 2538 2926 2572
rect 2960 2538 2998 2572
rect 3032 2538 3070 2572
rect 3104 2538 3142 2572
rect 3176 2538 3214 2572
rect 3248 2538 3286 2572
rect 3320 2538 3358 2572
rect 3392 2538 3430 2572
rect 3464 2538 3502 2572
rect 3536 2538 3574 2572
rect 3608 2538 3646 2572
rect 3680 2538 3718 2572
rect 3752 2538 3790 2572
rect 3824 2538 3862 2572
rect 3896 2538 3934 2572
rect 3968 2538 4006 2572
rect 4040 2538 4083 2572
rect 2091 2532 4083 2538
rect -4139 2465 -4093 2500
rect -4139 2431 -4133 2465
rect -4099 2431 -4093 2465
rect -4139 2393 -4093 2431
rect -4139 2359 -4133 2393
rect -4099 2359 -4093 2393
rect -4139 2321 -4093 2359
rect -4139 2287 -4133 2321
rect -4099 2287 -4093 2321
rect -4139 2249 -4093 2287
rect -4139 2215 -4133 2249
rect -4099 2215 -4093 2249
rect -4139 2177 -4093 2215
rect -4139 2143 -4133 2177
rect -4099 2143 -4093 2177
rect -4139 2105 -4093 2143
rect -4139 2071 -4133 2105
rect -4099 2071 -4093 2105
rect -4139 2033 -4093 2071
rect -4139 1999 -4133 2033
rect -4099 1999 -4093 2033
rect -4139 1961 -4093 1999
rect -4139 1927 -4133 1961
rect -4099 1927 -4093 1961
rect -4139 1889 -4093 1927
rect -4139 1855 -4133 1889
rect -4099 1855 -4093 1889
rect -4139 1817 -4093 1855
rect -4139 1783 -4133 1817
rect -4099 1783 -4093 1817
rect -4139 1745 -4093 1783
rect -4139 1711 -4133 1745
rect -4099 1711 -4093 1745
rect -4139 1673 -4093 1711
rect -4139 1639 -4133 1673
rect -4099 1639 -4093 1673
rect -4139 1601 -4093 1639
rect -4139 1567 -4133 1601
rect -4099 1567 -4093 1601
rect -4139 1529 -4093 1567
rect -4139 1495 -4133 1529
rect -4099 1495 -4093 1529
rect -4139 1457 -4093 1495
rect -4139 1423 -4133 1457
rect -4099 1423 -4093 1457
rect -4139 1385 -4093 1423
rect -4139 1351 -4133 1385
rect -4099 1351 -4093 1385
rect -4139 1313 -4093 1351
rect -4139 1279 -4133 1313
rect -4099 1279 -4093 1313
rect -4139 1241 -4093 1279
rect -4139 1207 -4133 1241
rect -4099 1207 -4093 1241
rect -4139 1169 -4093 1207
rect -4139 1135 -4133 1169
rect -4099 1135 -4093 1169
rect -4139 1097 -4093 1135
rect -4139 1063 -4133 1097
rect -4099 1063 -4093 1097
rect -4139 1025 -4093 1063
rect -4139 991 -4133 1025
rect -4099 991 -4093 1025
rect -4139 953 -4093 991
rect -4139 919 -4133 953
rect -4099 919 -4093 953
rect -4139 881 -4093 919
rect -4139 847 -4133 881
rect -4099 847 -4093 881
rect -4139 809 -4093 847
rect -4139 775 -4133 809
rect -4099 775 -4093 809
rect -4139 737 -4093 775
rect -4139 703 -4133 737
rect -4099 703 -4093 737
rect -4139 665 -4093 703
rect -4139 631 -4133 665
rect -4099 631 -4093 665
rect -4139 593 -4093 631
rect -4139 559 -4133 593
rect -4099 559 -4093 593
rect -4139 521 -4093 559
rect -4139 487 -4133 521
rect -4099 487 -4093 521
rect -4139 449 -4093 487
rect -4139 415 -4133 449
rect -4099 415 -4093 449
rect -4139 377 -4093 415
rect -4139 343 -4133 377
rect -4099 343 -4093 377
rect -4139 305 -4093 343
rect -4139 271 -4133 305
rect -4099 271 -4093 305
rect -4139 233 -4093 271
rect -4139 199 -4133 233
rect -4099 199 -4093 233
rect -4139 161 -4093 199
rect -4139 127 -4133 161
rect -4099 127 -4093 161
rect -4139 89 -4093 127
rect -4139 55 -4133 89
rect -4099 55 -4093 89
rect -4139 17 -4093 55
rect -4139 -17 -4133 17
rect -4099 -17 -4093 17
rect -4139 -55 -4093 -17
rect -4139 -89 -4133 -55
rect -4099 -89 -4093 -55
rect -4139 -127 -4093 -89
rect -4139 -161 -4133 -127
rect -4099 -161 -4093 -127
rect -4139 -199 -4093 -161
rect -4139 -233 -4133 -199
rect -4099 -233 -4093 -199
rect -4139 -271 -4093 -233
rect -4139 -305 -4133 -271
rect -4099 -305 -4093 -271
rect -4139 -343 -4093 -305
rect -4139 -377 -4133 -343
rect -4099 -377 -4093 -343
rect -4139 -415 -4093 -377
rect -4139 -449 -4133 -415
rect -4099 -449 -4093 -415
rect -4139 -487 -4093 -449
rect -4139 -521 -4133 -487
rect -4099 -521 -4093 -487
rect -4139 -559 -4093 -521
rect -4139 -593 -4133 -559
rect -4099 -593 -4093 -559
rect -4139 -631 -4093 -593
rect -4139 -665 -4133 -631
rect -4099 -665 -4093 -631
rect -4139 -703 -4093 -665
rect -4139 -737 -4133 -703
rect -4099 -737 -4093 -703
rect -4139 -775 -4093 -737
rect -4139 -809 -4133 -775
rect -4099 -809 -4093 -775
rect -4139 -847 -4093 -809
rect -4139 -881 -4133 -847
rect -4099 -881 -4093 -847
rect -4139 -919 -4093 -881
rect -4139 -953 -4133 -919
rect -4099 -953 -4093 -919
rect -4139 -991 -4093 -953
rect -4139 -1025 -4133 -991
rect -4099 -1025 -4093 -991
rect -4139 -1063 -4093 -1025
rect -4139 -1097 -4133 -1063
rect -4099 -1097 -4093 -1063
rect -4139 -1135 -4093 -1097
rect -4139 -1169 -4133 -1135
rect -4099 -1169 -4093 -1135
rect -4139 -1207 -4093 -1169
rect -4139 -1241 -4133 -1207
rect -4099 -1241 -4093 -1207
rect -4139 -1279 -4093 -1241
rect -4139 -1313 -4133 -1279
rect -4099 -1313 -4093 -1279
rect -4139 -1351 -4093 -1313
rect -4139 -1385 -4133 -1351
rect -4099 -1385 -4093 -1351
rect -4139 -1423 -4093 -1385
rect -4139 -1457 -4133 -1423
rect -4099 -1457 -4093 -1423
rect -4139 -1495 -4093 -1457
rect -4139 -1529 -4133 -1495
rect -4099 -1529 -4093 -1495
rect -4139 -1567 -4093 -1529
rect -4139 -1601 -4133 -1567
rect -4099 -1601 -4093 -1567
rect -4139 -1639 -4093 -1601
rect -4139 -1673 -4133 -1639
rect -4099 -1673 -4093 -1639
rect -4139 -1711 -4093 -1673
rect -4139 -1745 -4133 -1711
rect -4099 -1745 -4093 -1711
rect -4139 -1783 -4093 -1745
rect -4139 -1817 -4133 -1783
rect -4099 -1817 -4093 -1783
rect -4139 -1855 -4093 -1817
rect -4139 -1889 -4133 -1855
rect -4099 -1889 -4093 -1855
rect -4139 -1927 -4093 -1889
rect -4139 -1961 -4133 -1927
rect -4099 -1961 -4093 -1927
rect -4139 -1999 -4093 -1961
rect -4139 -2033 -4133 -1999
rect -4099 -2033 -4093 -1999
rect -4139 -2071 -4093 -2033
rect -4139 -2105 -4133 -2071
rect -4099 -2105 -4093 -2071
rect -4139 -2143 -4093 -2105
rect -4139 -2177 -4133 -2143
rect -4099 -2177 -4093 -2143
rect -4139 -2215 -4093 -2177
rect -4139 -2249 -4133 -2215
rect -4099 -2249 -4093 -2215
rect -4139 -2287 -4093 -2249
rect -4139 -2321 -4133 -2287
rect -4099 -2321 -4093 -2287
rect -4139 -2359 -4093 -2321
rect -4139 -2393 -4133 -2359
rect -4099 -2393 -4093 -2359
rect -4139 -2431 -4093 -2393
rect -4139 -2465 -4133 -2431
rect -4099 -2465 -4093 -2431
rect -4139 -2500 -4093 -2465
rect -2081 2465 -2035 2500
rect -2081 2431 -2075 2465
rect -2041 2431 -2035 2465
rect -2081 2393 -2035 2431
rect -2081 2359 -2075 2393
rect -2041 2359 -2035 2393
rect -2081 2321 -2035 2359
rect -2081 2287 -2075 2321
rect -2041 2287 -2035 2321
rect -2081 2249 -2035 2287
rect -2081 2215 -2075 2249
rect -2041 2215 -2035 2249
rect -2081 2177 -2035 2215
rect -2081 2143 -2075 2177
rect -2041 2143 -2035 2177
rect -2081 2105 -2035 2143
rect -2081 2071 -2075 2105
rect -2041 2071 -2035 2105
rect -2081 2033 -2035 2071
rect -2081 1999 -2075 2033
rect -2041 1999 -2035 2033
rect -2081 1961 -2035 1999
rect -2081 1927 -2075 1961
rect -2041 1927 -2035 1961
rect -2081 1889 -2035 1927
rect -2081 1855 -2075 1889
rect -2041 1855 -2035 1889
rect -2081 1817 -2035 1855
rect -2081 1783 -2075 1817
rect -2041 1783 -2035 1817
rect -2081 1745 -2035 1783
rect -2081 1711 -2075 1745
rect -2041 1711 -2035 1745
rect -2081 1673 -2035 1711
rect -2081 1639 -2075 1673
rect -2041 1639 -2035 1673
rect -2081 1601 -2035 1639
rect -2081 1567 -2075 1601
rect -2041 1567 -2035 1601
rect -2081 1529 -2035 1567
rect -2081 1495 -2075 1529
rect -2041 1495 -2035 1529
rect -2081 1457 -2035 1495
rect -2081 1423 -2075 1457
rect -2041 1423 -2035 1457
rect -2081 1385 -2035 1423
rect -2081 1351 -2075 1385
rect -2041 1351 -2035 1385
rect -2081 1313 -2035 1351
rect -2081 1279 -2075 1313
rect -2041 1279 -2035 1313
rect -2081 1241 -2035 1279
rect -2081 1207 -2075 1241
rect -2041 1207 -2035 1241
rect -2081 1169 -2035 1207
rect -2081 1135 -2075 1169
rect -2041 1135 -2035 1169
rect -2081 1097 -2035 1135
rect -2081 1063 -2075 1097
rect -2041 1063 -2035 1097
rect -2081 1025 -2035 1063
rect -2081 991 -2075 1025
rect -2041 991 -2035 1025
rect -2081 953 -2035 991
rect -2081 919 -2075 953
rect -2041 919 -2035 953
rect -2081 881 -2035 919
rect -2081 847 -2075 881
rect -2041 847 -2035 881
rect -2081 809 -2035 847
rect -2081 775 -2075 809
rect -2041 775 -2035 809
rect -2081 737 -2035 775
rect -2081 703 -2075 737
rect -2041 703 -2035 737
rect -2081 665 -2035 703
rect -2081 631 -2075 665
rect -2041 631 -2035 665
rect -2081 593 -2035 631
rect -2081 559 -2075 593
rect -2041 559 -2035 593
rect -2081 521 -2035 559
rect -2081 487 -2075 521
rect -2041 487 -2035 521
rect -2081 449 -2035 487
rect -2081 415 -2075 449
rect -2041 415 -2035 449
rect -2081 377 -2035 415
rect -2081 343 -2075 377
rect -2041 343 -2035 377
rect -2081 305 -2035 343
rect -2081 271 -2075 305
rect -2041 271 -2035 305
rect -2081 233 -2035 271
rect -2081 199 -2075 233
rect -2041 199 -2035 233
rect -2081 161 -2035 199
rect -2081 127 -2075 161
rect -2041 127 -2035 161
rect -2081 89 -2035 127
rect -2081 55 -2075 89
rect -2041 55 -2035 89
rect -2081 17 -2035 55
rect -2081 -17 -2075 17
rect -2041 -17 -2035 17
rect -2081 -55 -2035 -17
rect -2081 -89 -2075 -55
rect -2041 -89 -2035 -55
rect -2081 -127 -2035 -89
rect -2081 -161 -2075 -127
rect -2041 -161 -2035 -127
rect -2081 -199 -2035 -161
rect -2081 -233 -2075 -199
rect -2041 -233 -2035 -199
rect -2081 -271 -2035 -233
rect -2081 -305 -2075 -271
rect -2041 -305 -2035 -271
rect -2081 -343 -2035 -305
rect -2081 -377 -2075 -343
rect -2041 -377 -2035 -343
rect -2081 -415 -2035 -377
rect -2081 -449 -2075 -415
rect -2041 -449 -2035 -415
rect -2081 -487 -2035 -449
rect -2081 -521 -2075 -487
rect -2041 -521 -2035 -487
rect -2081 -559 -2035 -521
rect -2081 -593 -2075 -559
rect -2041 -593 -2035 -559
rect -2081 -631 -2035 -593
rect -2081 -665 -2075 -631
rect -2041 -665 -2035 -631
rect -2081 -703 -2035 -665
rect -2081 -737 -2075 -703
rect -2041 -737 -2035 -703
rect -2081 -775 -2035 -737
rect -2081 -809 -2075 -775
rect -2041 -809 -2035 -775
rect -2081 -847 -2035 -809
rect -2081 -881 -2075 -847
rect -2041 -881 -2035 -847
rect -2081 -919 -2035 -881
rect -2081 -953 -2075 -919
rect -2041 -953 -2035 -919
rect -2081 -991 -2035 -953
rect -2081 -1025 -2075 -991
rect -2041 -1025 -2035 -991
rect -2081 -1063 -2035 -1025
rect -2081 -1097 -2075 -1063
rect -2041 -1097 -2035 -1063
rect -2081 -1135 -2035 -1097
rect -2081 -1169 -2075 -1135
rect -2041 -1169 -2035 -1135
rect -2081 -1207 -2035 -1169
rect -2081 -1241 -2075 -1207
rect -2041 -1241 -2035 -1207
rect -2081 -1279 -2035 -1241
rect -2081 -1313 -2075 -1279
rect -2041 -1313 -2035 -1279
rect -2081 -1351 -2035 -1313
rect -2081 -1385 -2075 -1351
rect -2041 -1385 -2035 -1351
rect -2081 -1423 -2035 -1385
rect -2081 -1457 -2075 -1423
rect -2041 -1457 -2035 -1423
rect -2081 -1495 -2035 -1457
rect -2081 -1529 -2075 -1495
rect -2041 -1529 -2035 -1495
rect -2081 -1567 -2035 -1529
rect -2081 -1601 -2075 -1567
rect -2041 -1601 -2035 -1567
rect -2081 -1639 -2035 -1601
rect -2081 -1673 -2075 -1639
rect -2041 -1673 -2035 -1639
rect -2081 -1711 -2035 -1673
rect -2081 -1745 -2075 -1711
rect -2041 -1745 -2035 -1711
rect -2081 -1783 -2035 -1745
rect -2081 -1817 -2075 -1783
rect -2041 -1817 -2035 -1783
rect -2081 -1855 -2035 -1817
rect -2081 -1889 -2075 -1855
rect -2041 -1889 -2035 -1855
rect -2081 -1927 -2035 -1889
rect -2081 -1961 -2075 -1927
rect -2041 -1961 -2035 -1927
rect -2081 -1999 -2035 -1961
rect -2081 -2033 -2075 -1999
rect -2041 -2033 -2035 -1999
rect -2081 -2071 -2035 -2033
rect -2081 -2105 -2075 -2071
rect -2041 -2105 -2035 -2071
rect -2081 -2143 -2035 -2105
rect -2081 -2177 -2075 -2143
rect -2041 -2177 -2035 -2143
rect -2081 -2215 -2035 -2177
rect -2081 -2249 -2075 -2215
rect -2041 -2249 -2035 -2215
rect -2081 -2287 -2035 -2249
rect -2081 -2321 -2075 -2287
rect -2041 -2321 -2035 -2287
rect -2081 -2359 -2035 -2321
rect -2081 -2393 -2075 -2359
rect -2041 -2393 -2035 -2359
rect -2081 -2431 -2035 -2393
rect -2081 -2465 -2075 -2431
rect -2041 -2465 -2035 -2431
rect -2081 -2500 -2035 -2465
rect -23 2465 23 2500
rect -23 2431 -17 2465
rect 17 2431 23 2465
rect -23 2393 23 2431
rect -23 2359 -17 2393
rect 17 2359 23 2393
rect -23 2321 23 2359
rect -23 2287 -17 2321
rect 17 2287 23 2321
rect -23 2249 23 2287
rect -23 2215 -17 2249
rect 17 2215 23 2249
rect -23 2177 23 2215
rect -23 2143 -17 2177
rect 17 2143 23 2177
rect -23 2105 23 2143
rect -23 2071 -17 2105
rect 17 2071 23 2105
rect -23 2033 23 2071
rect -23 1999 -17 2033
rect 17 1999 23 2033
rect -23 1961 23 1999
rect -23 1927 -17 1961
rect 17 1927 23 1961
rect -23 1889 23 1927
rect -23 1855 -17 1889
rect 17 1855 23 1889
rect -23 1817 23 1855
rect -23 1783 -17 1817
rect 17 1783 23 1817
rect -23 1745 23 1783
rect -23 1711 -17 1745
rect 17 1711 23 1745
rect -23 1673 23 1711
rect -23 1639 -17 1673
rect 17 1639 23 1673
rect -23 1601 23 1639
rect -23 1567 -17 1601
rect 17 1567 23 1601
rect -23 1529 23 1567
rect -23 1495 -17 1529
rect 17 1495 23 1529
rect -23 1457 23 1495
rect -23 1423 -17 1457
rect 17 1423 23 1457
rect -23 1385 23 1423
rect -23 1351 -17 1385
rect 17 1351 23 1385
rect -23 1313 23 1351
rect -23 1279 -17 1313
rect 17 1279 23 1313
rect -23 1241 23 1279
rect -23 1207 -17 1241
rect 17 1207 23 1241
rect -23 1169 23 1207
rect -23 1135 -17 1169
rect 17 1135 23 1169
rect -23 1097 23 1135
rect -23 1063 -17 1097
rect 17 1063 23 1097
rect -23 1025 23 1063
rect -23 991 -17 1025
rect 17 991 23 1025
rect -23 953 23 991
rect -23 919 -17 953
rect 17 919 23 953
rect -23 881 23 919
rect -23 847 -17 881
rect 17 847 23 881
rect -23 809 23 847
rect -23 775 -17 809
rect 17 775 23 809
rect -23 737 23 775
rect -23 703 -17 737
rect 17 703 23 737
rect -23 665 23 703
rect -23 631 -17 665
rect 17 631 23 665
rect -23 593 23 631
rect -23 559 -17 593
rect 17 559 23 593
rect -23 521 23 559
rect -23 487 -17 521
rect 17 487 23 521
rect -23 449 23 487
rect -23 415 -17 449
rect 17 415 23 449
rect -23 377 23 415
rect -23 343 -17 377
rect 17 343 23 377
rect -23 305 23 343
rect -23 271 -17 305
rect 17 271 23 305
rect -23 233 23 271
rect -23 199 -17 233
rect 17 199 23 233
rect -23 161 23 199
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -199 23 -161
rect -23 -233 -17 -199
rect 17 -233 23 -199
rect -23 -271 23 -233
rect -23 -305 -17 -271
rect 17 -305 23 -271
rect -23 -343 23 -305
rect -23 -377 -17 -343
rect 17 -377 23 -343
rect -23 -415 23 -377
rect -23 -449 -17 -415
rect 17 -449 23 -415
rect -23 -487 23 -449
rect -23 -521 -17 -487
rect 17 -521 23 -487
rect -23 -559 23 -521
rect -23 -593 -17 -559
rect 17 -593 23 -559
rect -23 -631 23 -593
rect -23 -665 -17 -631
rect 17 -665 23 -631
rect -23 -703 23 -665
rect -23 -737 -17 -703
rect 17 -737 23 -703
rect -23 -775 23 -737
rect -23 -809 -17 -775
rect 17 -809 23 -775
rect -23 -847 23 -809
rect -23 -881 -17 -847
rect 17 -881 23 -847
rect -23 -919 23 -881
rect -23 -953 -17 -919
rect 17 -953 23 -919
rect -23 -991 23 -953
rect -23 -1025 -17 -991
rect 17 -1025 23 -991
rect -23 -1063 23 -1025
rect -23 -1097 -17 -1063
rect 17 -1097 23 -1063
rect -23 -1135 23 -1097
rect -23 -1169 -17 -1135
rect 17 -1169 23 -1135
rect -23 -1207 23 -1169
rect -23 -1241 -17 -1207
rect 17 -1241 23 -1207
rect -23 -1279 23 -1241
rect -23 -1313 -17 -1279
rect 17 -1313 23 -1279
rect -23 -1351 23 -1313
rect -23 -1385 -17 -1351
rect 17 -1385 23 -1351
rect -23 -1423 23 -1385
rect -23 -1457 -17 -1423
rect 17 -1457 23 -1423
rect -23 -1495 23 -1457
rect -23 -1529 -17 -1495
rect 17 -1529 23 -1495
rect -23 -1567 23 -1529
rect -23 -1601 -17 -1567
rect 17 -1601 23 -1567
rect -23 -1639 23 -1601
rect -23 -1673 -17 -1639
rect 17 -1673 23 -1639
rect -23 -1711 23 -1673
rect -23 -1745 -17 -1711
rect 17 -1745 23 -1711
rect -23 -1783 23 -1745
rect -23 -1817 -17 -1783
rect 17 -1817 23 -1783
rect -23 -1855 23 -1817
rect -23 -1889 -17 -1855
rect 17 -1889 23 -1855
rect -23 -1927 23 -1889
rect -23 -1961 -17 -1927
rect 17 -1961 23 -1927
rect -23 -1999 23 -1961
rect -23 -2033 -17 -1999
rect 17 -2033 23 -1999
rect -23 -2071 23 -2033
rect -23 -2105 -17 -2071
rect 17 -2105 23 -2071
rect -23 -2143 23 -2105
rect -23 -2177 -17 -2143
rect 17 -2177 23 -2143
rect -23 -2215 23 -2177
rect -23 -2249 -17 -2215
rect 17 -2249 23 -2215
rect -23 -2287 23 -2249
rect -23 -2321 -17 -2287
rect 17 -2321 23 -2287
rect -23 -2359 23 -2321
rect -23 -2393 -17 -2359
rect 17 -2393 23 -2359
rect -23 -2431 23 -2393
rect -23 -2465 -17 -2431
rect 17 -2465 23 -2431
rect -23 -2500 23 -2465
rect 2035 2465 2081 2500
rect 2035 2431 2041 2465
rect 2075 2431 2081 2465
rect 2035 2393 2081 2431
rect 2035 2359 2041 2393
rect 2075 2359 2081 2393
rect 2035 2321 2081 2359
rect 2035 2287 2041 2321
rect 2075 2287 2081 2321
rect 2035 2249 2081 2287
rect 2035 2215 2041 2249
rect 2075 2215 2081 2249
rect 2035 2177 2081 2215
rect 2035 2143 2041 2177
rect 2075 2143 2081 2177
rect 2035 2105 2081 2143
rect 2035 2071 2041 2105
rect 2075 2071 2081 2105
rect 2035 2033 2081 2071
rect 2035 1999 2041 2033
rect 2075 1999 2081 2033
rect 2035 1961 2081 1999
rect 2035 1927 2041 1961
rect 2075 1927 2081 1961
rect 2035 1889 2081 1927
rect 2035 1855 2041 1889
rect 2075 1855 2081 1889
rect 2035 1817 2081 1855
rect 2035 1783 2041 1817
rect 2075 1783 2081 1817
rect 2035 1745 2081 1783
rect 2035 1711 2041 1745
rect 2075 1711 2081 1745
rect 2035 1673 2081 1711
rect 2035 1639 2041 1673
rect 2075 1639 2081 1673
rect 2035 1601 2081 1639
rect 2035 1567 2041 1601
rect 2075 1567 2081 1601
rect 2035 1529 2081 1567
rect 2035 1495 2041 1529
rect 2075 1495 2081 1529
rect 2035 1457 2081 1495
rect 2035 1423 2041 1457
rect 2075 1423 2081 1457
rect 2035 1385 2081 1423
rect 2035 1351 2041 1385
rect 2075 1351 2081 1385
rect 2035 1313 2081 1351
rect 2035 1279 2041 1313
rect 2075 1279 2081 1313
rect 2035 1241 2081 1279
rect 2035 1207 2041 1241
rect 2075 1207 2081 1241
rect 2035 1169 2081 1207
rect 2035 1135 2041 1169
rect 2075 1135 2081 1169
rect 2035 1097 2081 1135
rect 2035 1063 2041 1097
rect 2075 1063 2081 1097
rect 2035 1025 2081 1063
rect 2035 991 2041 1025
rect 2075 991 2081 1025
rect 2035 953 2081 991
rect 2035 919 2041 953
rect 2075 919 2081 953
rect 2035 881 2081 919
rect 2035 847 2041 881
rect 2075 847 2081 881
rect 2035 809 2081 847
rect 2035 775 2041 809
rect 2075 775 2081 809
rect 2035 737 2081 775
rect 2035 703 2041 737
rect 2075 703 2081 737
rect 2035 665 2081 703
rect 2035 631 2041 665
rect 2075 631 2081 665
rect 2035 593 2081 631
rect 2035 559 2041 593
rect 2075 559 2081 593
rect 2035 521 2081 559
rect 2035 487 2041 521
rect 2075 487 2081 521
rect 2035 449 2081 487
rect 2035 415 2041 449
rect 2075 415 2081 449
rect 2035 377 2081 415
rect 2035 343 2041 377
rect 2075 343 2081 377
rect 2035 305 2081 343
rect 2035 271 2041 305
rect 2075 271 2081 305
rect 2035 233 2081 271
rect 2035 199 2041 233
rect 2075 199 2081 233
rect 2035 161 2081 199
rect 2035 127 2041 161
rect 2075 127 2081 161
rect 2035 89 2081 127
rect 2035 55 2041 89
rect 2075 55 2081 89
rect 2035 17 2081 55
rect 2035 -17 2041 17
rect 2075 -17 2081 17
rect 2035 -55 2081 -17
rect 2035 -89 2041 -55
rect 2075 -89 2081 -55
rect 2035 -127 2081 -89
rect 2035 -161 2041 -127
rect 2075 -161 2081 -127
rect 2035 -199 2081 -161
rect 2035 -233 2041 -199
rect 2075 -233 2081 -199
rect 2035 -271 2081 -233
rect 2035 -305 2041 -271
rect 2075 -305 2081 -271
rect 2035 -343 2081 -305
rect 2035 -377 2041 -343
rect 2075 -377 2081 -343
rect 2035 -415 2081 -377
rect 2035 -449 2041 -415
rect 2075 -449 2081 -415
rect 2035 -487 2081 -449
rect 2035 -521 2041 -487
rect 2075 -521 2081 -487
rect 2035 -559 2081 -521
rect 2035 -593 2041 -559
rect 2075 -593 2081 -559
rect 2035 -631 2081 -593
rect 2035 -665 2041 -631
rect 2075 -665 2081 -631
rect 2035 -703 2081 -665
rect 2035 -737 2041 -703
rect 2075 -737 2081 -703
rect 2035 -775 2081 -737
rect 2035 -809 2041 -775
rect 2075 -809 2081 -775
rect 2035 -847 2081 -809
rect 2035 -881 2041 -847
rect 2075 -881 2081 -847
rect 2035 -919 2081 -881
rect 2035 -953 2041 -919
rect 2075 -953 2081 -919
rect 2035 -991 2081 -953
rect 2035 -1025 2041 -991
rect 2075 -1025 2081 -991
rect 2035 -1063 2081 -1025
rect 2035 -1097 2041 -1063
rect 2075 -1097 2081 -1063
rect 2035 -1135 2081 -1097
rect 2035 -1169 2041 -1135
rect 2075 -1169 2081 -1135
rect 2035 -1207 2081 -1169
rect 2035 -1241 2041 -1207
rect 2075 -1241 2081 -1207
rect 2035 -1279 2081 -1241
rect 2035 -1313 2041 -1279
rect 2075 -1313 2081 -1279
rect 2035 -1351 2081 -1313
rect 2035 -1385 2041 -1351
rect 2075 -1385 2081 -1351
rect 2035 -1423 2081 -1385
rect 2035 -1457 2041 -1423
rect 2075 -1457 2081 -1423
rect 2035 -1495 2081 -1457
rect 2035 -1529 2041 -1495
rect 2075 -1529 2081 -1495
rect 2035 -1567 2081 -1529
rect 2035 -1601 2041 -1567
rect 2075 -1601 2081 -1567
rect 2035 -1639 2081 -1601
rect 2035 -1673 2041 -1639
rect 2075 -1673 2081 -1639
rect 2035 -1711 2081 -1673
rect 2035 -1745 2041 -1711
rect 2075 -1745 2081 -1711
rect 2035 -1783 2081 -1745
rect 2035 -1817 2041 -1783
rect 2075 -1817 2081 -1783
rect 2035 -1855 2081 -1817
rect 2035 -1889 2041 -1855
rect 2075 -1889 2081 -1855
rect 2035 -1927 2081 -1889
rect 2035 -1961 2041 -1927
rect 2075 -1961 2081 -1927
rect 2035 -1999 2081 -1961
rect 2035 -2033 2041 -1999
rect 2075 -2033 2081 -1999
rect 2035 -2071 2081 -2033
rect 2035 -2105 2041 -2071
rect 2075 -2105 2081 -2071
rect 2035 -2143 2081 -2105
rect 2035 -2177 2041 -2143
rect 2075 -2177 2081 -2143
rect 2035 -2215 2081 -2177
rect 2035 -2249 2041 -2215
rect 2075 -2249 2081 -2215
rect 2035 -2287 2081 -2249
rect 2035 -2321 2041 -2287
rect 2075 -2321 2081 -2287
rect 2035 -2359 2081 -2321
rect 2035 -2393 2041 -2359
rect 2075 -2393 2081 -2359
rect 2035 -2431 2081 -2393
rect 2035 -2465 2041 -2431
rect 2075 -2465 2081 -2431
rect 2035 -2500 2081 -2465
rect 4093 2465 4139 2500
rect 4093 2431 4099 2465
rect 4133 2431 4139 2465
rect 4093 2393 4139 2431
rect 4093 2359 4099 2393
rect 4133 2359 4139 2393
rect 4093 2321 4139 2359
rect 4093 2287 4099 2321
rect 4133 2287 4139 2321
rect 4093 2249 4139 2287
rect 4093 2215 4099 2249
rect 4133 2215 4139 2249
rect 4093 2177 4139 2215
rect 4093 2143 4099 2177
rect 4133 2143 4139 2177
rect 4093 2105 4139 2143
rect 4093 2071 4099 2105
rect 4133 2071 4139 2105
rect 4093 2033 4139 2071
rect 4093 1999 4099 2033
rect 4133 1999 4139 2033
rect 4093 1961 4139 1999
rect 4093 1927 4099 1961
rect 4133 1927 4139 1961
rect 4093 1889 4139 1927
rect 4093 1855 4099 1889
rect 4133 1855 4139 1889
rect 4093 1817 4139 1855
rect 4093 1783 4099 1817
rect 4133 1783 4139 1817
rect 4093 1745 4139 1783
rect 4093 1711 4099 1745
rect 4133 1711 4139 1745
rect 4093 1673 4139 1711
rect 4093 1639 4099 1673
rect 4133 1639 4139 1673
rect 4093 1601 4139 1639
rect 4093 1567 4099 1601
rect 4133 1567 4139 1601
rect 4093 1529 4139 1567
rect 4093 1495 4099 1529
rect 4133 1495 4139 1529
rect 4093 1457 4139 1495
rect 4093 1423 4099 1457
rect 4133 1423 4139 1457
rect 4093 1385 4139 1423
rect 4093 1351 4099 1385
rect 4133 1351 4139 1385
rect 4093 1313 4139 1351
rect 4093 1279 4099 1313
rect 4133 1279 4139 1313
rect 4093 1241 4139 1279
rect 4093 1207 4099 1241
rect 4133 1207 4139 1241
rect 4093 1169 4139 1207
rect 4093 1135 4099 1169
rect 4133 1135 4139 1169
rect 4093 1097 4139 1135
rect 4093 1063 4099 1097
rect 4133 1063 4139 1097
rect 4093 1025 4139 1063
rect 4093 991 4099 1025
rect 4133 991 4139 1025
rect 4093 953 4139 991
rect 4093 919 4099 953
rect 4133 919 4139 953
rect 4093 881 4139 919
rect 4093 847 4099 881
rect 4133 847 4139 881
rect 4093 809 4139 847
rect 4093 775 4099 809
rect 4133 775 4139 809
rect 4093 737 4139 775
rect 4093 703 4099 737
rect 4133 703 4139 737
rect 4093 665 4139 703
rect 4093 631 4099 665
rect 4133 631 4139 665
rect 4093 593 4139 631
rect 4093 559 4099 593
rect 4133 559 4139 593
rect 4093 521 4139 559
rect 4093 487 4099 521
rect 4133 487 4139 521
rect 4093 449 4139 487
rect 4093 415 4099 449
rect 4133 415 4139 449
rect 4093 377 4139 415
rect 4093 343 4099 377
rect 4133 343 4139 377
rect 4093 305 4139 343
rect 4093 271 4099 305
rect 4133 271 4139 305
rect 4093 233 4139 271
rect 4093 199 4099 233
rect 4133 199 4139 233
rect 4093 161 4139 199
rect 4093 127 4099 161
rect 4133 127 4139 161
rect 4093 89 4139 127
rect 4093 55 4099 89
rect 4133 55 4139 89
rect 4093 17 4139 55
rect 4093 -17 4099 17
rect 4133 -17 4139 17
rect 4093 -55 4139 -17
rect 4093 -89 4099 -55
rect 4133 -89 4139 -55
rect 4093 -127 4139 -89
rect 4093 -161 4099 -127
rect 4133 -161 4139 -127
rect 4093 -199 4139 -161
rect 4093 -233 4099 -199
rect 4133 -233 4139 -199
rect 4093 -271 4139 -233
rect 4093 -305 4099 -271
rect 4133 -305 4139 -271
rect 4093 -343 4139 -305
rect 4093 -377 4099 -343
rect 4133 -377 4139 -343
rect 4093 -415 4139 -377
rect 4093 -449 4099 -415
rect 4133 -449 4139 -415
rect 4093 -487 4139 -449
rect 4093 -521 4099 -487
rect 4133 -521 4139 -487
rect 4093 -559 4139 -521
rect 4093 -593 4099 -559
rect 4133 -593 4139 -559
rect 4093 -631 4139 -593
rect 4093 -665 4099 -631
rect 4133 -665 4139 -631
rect 4093 -703 4139 -665
rect 4093 -737 4099 -703
rect 4133 -737 4139 -703
rect 4093 -775 4139 -737
rect 4093 -809 4099 -775
rect 4133 -809 4139 -775
rect 4093 -847 4139 -809
rect 4093 -881 4099 -847
rect 4133 -881 4139 -847
rect 4093 -919 4139 -881
rect 4093 -953 4099 -919
rect 4133 -953 4139 -919
rect 4093 -991 4139 -953
rect 4093 -1025 4099 -991
rect 4133 -1025 4139 -991
rect 4093 -1063 4139 -1025
rect 4093 -1097 4099 -1063
rect 4133 -1097 4139 -1063
rect 4093 -1135 4139 -1097
rect 4093 -1169 4099 -1135
rect 4133 -1169 4139 -1135
rect 4093 -1207 4139 -1169
rect 4093 -1241 4099 -1207
rect 4133 -1241 4139 -1207
rect 4093 -1279 4139 -1241
rect 4093 -1313 4099 -1279
rect 4133 -1313 4139 -1279
rect 4093 -1351 4139 -1313
rect 4093 -1385 4099 -1351
rect 4133 -1385 4139 -1351
rect 4093 -1423 4139 -1385
rect 4093 -1457 4099 -1423
rect 4133 -1457 4139 -1423
rect 4093 -1495 4139 -1457
rect 4093 -1529 4099 -1495
rect 4133 -1529 4139 -1495
rect 4093 -1567 4139 -1529
rect 4093 -1601 4099 -1567
rect 4133 -1601 4139 -1567
rect 4093 -1639 4139 -1601
rect 4093 -1673 4099 -1639
rect 4133 -1673 4139 -1639
rect 4093 -1711 4139 -1673
rect 4093 -1745 4099 -1711
rect 4133 -1745 4139 -1711
rect 4093 -1783 4139 -1745
rect 4093 -1817 4099 -1783
rect 4133 -1817 4139 -1783
rect 4093 -1855 4139 -1817
rect 4093 -1889 4099 -1855
rect 4133 -1889 4139 -1855
rect 4093 -1927 4139 -1889
rect 4093 -1961 4099 -1927
rect 4133 -1961 4139 -1927
rect 4093 -1999 4139 -1961
rect 4093 -2033 4099 -1999
rect 4133 -2033 4139 -1999
rect 4093 -2071 4139 -2033
rect 4093 -2105 4099 -2071
rect 4133 -2105 4139 -2071
rect 4093 -2143 4139 -2105
rect 4093 -2177 4099 -2143
rect 4133 -2177 4139 -2143
rect 4093 -2215 4139 -2177
rect 4093 -2249 4099 -2215
rect 4133 -2249 4139 -2215
rect 4093 -2287 4139 -2249
rect 4093 -2321 4099 -2287
rect 4133 -2321 4139 -2287
rect 4093 -2359 4139 -2321
rect 4093 -2393 4099 -2359
rect 4133 -2393 4139 -2359
rect 4093 -2431 4139 -2393
rect 4093 -2465 4099 -2431
rect 4133 -2465 4139 -2431
rect 4093 -2500 4139 -2465
rect -4083 -2538 -2091 -2532
rect -4083 -2572 -4040 -2538
rect -4006 -2572 -3968 -2538
rect -3934 -2572 -3896 -2538
rect -3862 -2572 -3824 -2538
rect -3790 -2572 -3752 -2538
rect -3718 -2572 -3680 -2538
rect -3646 -2572 -3608 -2538
rect -3574 -2572 -3536 -2538
rect -3502 -2572 -3464 -2538
rect -3430 -2572 -3392 -2538
rect -3358 -2572 -3320 -2538
rect -3286 -2572 -3248 -2538
rect -3214 -2572 -3176 -2538
rect -3142 -2572 -3104 -2538
rect -3070 -2572 -3032 -2538
rect -2998 -2572 -2960 -2538
rect -2926 -2572 -2888 -2538
rect -2854 -2572 -2816 -2538
rect -2782 -2572 -2744 -2538
rect -2710 -2572 -2672 -2538
rect -2638 -2572 -2600 -2538
rect -2566 -2572 -2528 -2538
rect -2494 -2572 -2456 -2538
rect -2422 -2572 -2384 -2538
rect -2350 -2572 -2312 -2538
rect -2278 -2572 -2240 -2538
rect -2206 -2572 -2168 -2538
rect -2134 -2572 -2091 -2538
rect -4083 -2578 -2091 -2572
rect -2025 -2538 -33 -2532
rect -2025 -2572 -1982 -2538
rect -1948 -2572 -1910 -2538
rect -1876 -2572 -1838 -2538
rect -1804 -2572 -1766 -2538
rect -1732 -2572 -1694 -2538
rect -1660 -2572 -1622 -2538
rect -1588 -2572 -1550 -2538
rect -1516 -2572 -1478 -2538
rect -1444 -2572 -1406 -2538
rect -1372 -2572 -1334 -2538
rect -1300 -2572 -1262 -2538
rect -1228 -2572 -1190 -2538
rect -1156 -2572 -1118 -2538
rect -1084 -2572 -1046 -2538
rect -1012 -2572 -974 -2538
rect -940 -2572 -902 -2538
rect -868 -2572 -830 -2538
rect -796 -2572 -758 -2538
rect -724 -2572 -686 -2538
rect -652 -2572 -614 -2538
rect -580 -2572 -542 -2538
rect -508 -2572 -470 -2538
rect -436 -2572 -398 -2538
rect -364 -2572 -326 -2538
rect -292 -2572 -254 -2538
rect -220 -2572 -182 -2538
rect -148 -2572 -110 -2538
rect -76 -2572 -33 -2538
rect -2025 -2578 -33 -2572
rect 33 -2538 2025 -2532
rect 33 -2572 76 -2538
rect 110 -2572 148 -2538
rect 182 -2572 220 -2538
rect 254 -2572 292 -2538
rect 326 -2572 364 -2538
rect 398 -2572 436 -2538
rect 470 -2572 508 -2538
rect 542 -2572 580 -2538
rect 614 -2572 652 -2538
rect 686 -2572 724 -2538
rect 758 -2572 796 -2538
rect 830 -2572 868 -2538
rect 902 -2572 940 -2538
rect 974 -2572 1012 -2538
rect 1046 -2572 1084 -2538
rect 1118 -2572 1156 -2538
rect 1190 -2572 1228 -2538
rect 1262 -2572 1300 -2538
rect 1334 -2572 1372 -2538
rect 1406 -2572 1444 -2538
rect 1478 -2572 1516 -2538
rect 1550 -2572 1588 -2538
rect 1622 -2572 1660 -2538
rect 1694 -2572 1732 -2538
rect 1766 -2572 1804 -2538
rect 1838 -2572 1876 -2538
rect 1910 -2572 1948 -2538
rect 1982 -2572 2025 -2538
rect 33 -2578 2025 -2572
rect 2091 -2538 4083 -2532
rect 2091 -2572 2134 -2538
rect 2168 -2572 2206 -2538
rect 2240 -2572 2278 -2538
rect 2312 -2572 2350 -2538
rect 2384 -2572 2422 -2538
rect 2456 -2572 2494 -2538
rect 2528 -2572 2566 -2538
rect 2600 -2572 2638 -2538
rect 2672 -2572 2710 -2538
rect 2744 -2572 2782 -2538
rect 2816 -2572 2854 -2538
rect 2888 -2572 2926 -2538
rect 2960 -2572 2998 -2538
rect 3032 -2572 3070 -2538
rect 3104 -2572 3142 -2538
rect 3176 -2572 3214 -2538
rect 3248 -2572 3286 -2538
rect 3320 -2572 3358 -2538
rect 3392 -2572 3430 -2538
rect 3464 -2572 3502 -2538
rect 3536 -2572 3574 -2538
rect 3608 -2572 3646 -2538
rect 3680 -2572 3718 -2538
rect 3752 -2572 3790 -2538
rect 3824 -2572 3862 -2538
rect 3896 -2572 3934 -2538
rect 3968 -2572 4006 -2538
rect 4040 -2572 4083 -2538
rect 2091 -2578 4083 -2572
<< properties >>
string FIXED_BBOX -4230 -2657 4230 2657
<< end >>
