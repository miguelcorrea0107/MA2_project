magic
tech sky130A
magscale 1 2
timestamp 1716644424
<< pwell >>
rect -1447 -2700 1447 2700
<< nmos >>
rect -1261 -2500 -1061 2500
rect -1003 -2500 -803 2500
rect -745 -2500 -545 2500
rect -487 -2500 -287 2500
rect -229 -2500 -29 2500
rect 29 -2500 229 2500
rect 287 -2500 487 2500
rect 545 -2500 745 2500
rect 803 -2500 1003 2500
rect 1061 -2500 1261 2500
<< ndiff >>
rect -1319 2465 -1261 2500
rect -1319 2431 -1307 2465
rect -1273 2431 -1261 2465
rect -1319 2397 -1261 2431
rect -1319 2363 -1307 2397
rect -1273 2363 -1261 2397
rect -1319 2329 -1261 2363
rect -1319 2295 -1307 2329
rect -1273 2295 -1261 2329
rect -1319 2261 -1261 2295
rect -1319 2227 -1307 2261
rect -1273 2227 -1261 2261
rect -1319 2193 -1261 2227
rect -1319 2159 -1307 2193
rect -1273 2159 -1261 2193
rect -1319 2125 -1261 2159
rect -1319 2091 -1307 2125
rect -1273 2091 -1261 2125
rect -1319 2057 -1261 2091
rect -1319 2023 -1307 2057
rect -1273 2023 -1261 2057
rect -1319 1989 -1261 2023
rect -1319 1955 -1307 1989
rect -1273 1955 -1261 1989
rect -1319 1921 -1261 1955
rect -1319 1887 -1307 1921
rect -1273 1887 -1261 1921
rect -1319 1853 -1261 1887
rect -1319 1819 -1307 1853
rect -1273 1819 -1261 1853
rect -1319 1785 -1261 1819
rect -1319 1751 -1307 1785
rect -1273 1751 -1261 1785
rect -1319 1717 -1261 1751
rect -1319 1683 -1307 1717
rect -1273 1683 -1261 1717
rect -1319 1649 -1261 1683
rect -1319 1615 -1307 1649
rect -1273 1615 -1261 1649
rect -1319 1581 -1261 1615
rect -1319 1547 -1307 1581
rect -1273 1547 -1261 1581
rect -1319 1513 -1261 1547
rect -1319 1479 -1307 1513
rect -1273 1479 -1261 1513
rect -1319 1445 -1261 1479
rect -1319 1411 -1307 1445
rect -1273 1411 -1261 1445
rect -1319 1377 -1261 1411
rect -1319 1343 -1307 1377
rect -1273 1343 -1261 1377
rect -1319 1309 -1261 1343
rect -1319 1275 -1307 1309
rect -1273 1275 -1261 1309
rect -1319 1241 -1261 1275
rect -1319 1207 -1307 1241
rect -1273 1207 -1261 1241
rect -1319 1173 -1261 1207
rect -1319 1139 -1307 1173
rect -1273 1139 -1261 1173
rect -1319 1105 -1261 1139
rect -1319 1071 -1307 1105
rect -1273 1071 -1261 1105
rect -1319 1037 -1261 1071
rect -1319 1003 -1307 1037
rect -1273 1003 -1261 1037
rect -1319 969 -1261 1003
rect -1319 935 -1307 969
rect -1273 935 -1261 969
rect -1319 901 -1261 935
rect -1319 867 -1307 901
rect -1273 867 -1261 901
rect -1319 833 -1261 867
rect -1319 799 -1307 833
rect -1273 799 -1261 833
rect -1319 765 -1261 799
rect -1319 731 -1307 765
rect -1273 731 -1261 765
rect -1319 697 -1261 731
rect -1319 663 -1307 697
rect -1273 663 -1261 697
rect -1319 629 -1261 663
rect -1319 595 -1307 629
rect -1273 595 -1261 629
rect -1319 561 -1261 595
rect -1319 527 -1307 561
rect -1273 527 -1261 561
rect -1319 493 -1261 527
rect -1319 459 -1307 493
rect -1273 459 -1261 493
rect -1319 425 -1261 459
rect -1319 391 -1307 425
rect -1273 391 -1261 425
rect -1319 357 -1261 391
rect -1319 323 -1307 357
rect -1273 323 -1261 357
rect -1319 289 -1261 323
rect -1319 255 -1307 289
rect -1273 255 -1261 289
rect -1319 221 -1261 255
rect -1319 187 -1307 221
rect -1273 187 -1261 221
rect -1319 153 -1261 187
rect -1319 119 -1307 153
rect -1273 119 -1261 153
rect -1319 85 -1261 119
rect -1319 51 -1307 85
rect -1273 51 -1261 85
rect -1319 17 -1261 51
rect -1319 -17 -1307 17
rect -1273 -17 -1261 17
rect -1319 -51 -1261 -17
rect -1319 -85 -1307 -51
rect -1273 -85 -1261 -51
rect -1319 -119 -1261 -85
rect -1319 -153 -1307 -119
rect -1273 -153 -1261 -119
rect -1319 -187 -1261 -153
rect -1319 -221 -1307 -187
rect -1273 -221 -1261 -187
rect -1319 -255 -1261 -221
rect -1319 -289 -1307 -255
rect -1273 -289 -1261 -255
rect -1319 -323 -1261 -289
rect -1319 -357 -1307 -323
rect -1273 -357 -1261 -323
rect -1319 -391 -1261 -357
rect -1319 -425 -1307 -391
rect -1273 -425 -1261 -391
rect -1319 -459 -1261 -425
rect -1319 -493 -1307 -459
rect -1273 -493 -1261 -459
rect -1319 -527 -1261 -493
rect -1319 -561 -1307 -527
rect -1273 -561 -1261 -527
rect -1319 -595 -1261 -561
rect -1319 -629 -1307 -595
rect -1273 -629 -1261 -595
rect -1319 -663 -1261 -629
rect -1319 -697 -1307 -663
rect -1273 -697 -1261 -663
rect -1319 -731 -1261 -697
rect -1319 -765 -1307 -731
rect -1273 -765 -1261 -731
rect -1319 -799 -1261 -765
rect -1319 -833 -1307 -799
rect -1273 -833 -1261 -799
rect -1319 -867 -1261 -833
rect -1319 -901 -1307 -867
rect -1273 -901 -1261 -867
rect -1319 -935 -1261 -901
rect -1319 -969 -1307 -935
rect -1273 -969 -1261 -935
rect -1319 -1003 -1261 -969
rect -1319 -1037 -1307 -1003
rect -1273 -1037 -1261 -1003
rect -1319 -1071 -1261 -1037
rect -1319 -1105 -1307 -1071
rect -1273 -1105 -1261 -1071
rect -1319 -1139 -1261 -1105
rect -1319 -1173 -1307 -1139
rect -1273 -1173 -1261 -1139
rect -1319 -1207 -1261 -1173
rect -1319 -1241 -1307 -1207
rect -1273 -1241 -1261 -1207
rect -1319 -1275 -1261 -1241
rect -1319 -1309 -1307 -1275
rect -1273 -1309 -1261 -1275
rect -1319 -1343 -1261 -1309
rect -1319 -1377 -1307 -1343
rect -1273 -1377 -1261 -1343
rect -1319 -1411 -1261 -1377
rect -1319 -1445 -1307 -1411
rect -1273 -1445 -1261 -1411
rect -1319 -1479 -1261 -1445
rect -1319 -1513 -1307 -1479
rect -1273 -1513 -1261 -1479
rect -1319 -1547 -1261 -1513
rect -1319 -1581 -1307 -1547
rect -1273 -1581 -1261 -1547
rect -1319 -1615 -1261 -1581
rect -1319 -1649 -1307 -1615
rect -1273 -1649 -1261 -1615
rect -1319 -1683 -1261 -1649
rect -1319 -1717 -1307 -1683
rect -1273 -1717 -1261 -1683
rect -1319 -1751 -1261 -1717
rect -1319 -1785 -1307 -1751
rect -1273 -1785 -1261 -1751
rect -1319 -1819 -1261 -1785
rect -1319 -1853 -1307 -1819
rect -1273 -1853 -1261 -1819
rect -1319 -1887 -1261 -1853
rect -1319 -1921 -1307 -1887
rect -1273 -1921 -1261 -1887
rect -1319 -1955 -1261 -1921
rect -1319 -1989 -1307 -1955
rect -1273 -1989 -1261 -1955
rect -1319 -2023 -1261 -1989
rect -1319 -2057 -1307 -2023
rect -1273 -2057 -1261 -2023
rect -1319 -2091 -1261 -2057
rect -1319 -2125 -1307 -2091
rect -1273 -2125 -1261 -2091
rect -1319 -2159 -1261 -2125
rect -1319 -2193 -1307 -2159
rect -1273 -2193 -1261 -2159
rect -1319 -2227 -1261 -2193
rect -1319 -2261 -1307 -2227
rect -1273 -2261 -1261 -2227
rect -1319 -2295 -1261 -2261
rect -1319 -2329 -1307 -2295
rect -1273 -2329 -1261 -2295
rect -1319 -2363 -1261 -2329
rect -1319 -2397 -1307 -2363
rect -1273 -2397 -1261 -2363
rect -1319 -2431 -1261 -2397
rect -1319 -2465 -1307 -2431
rect -1273 -2465 -1261 -2431
rect -1319 -2500 -1261 -2465
rect -1061 2465 -1003 2500
rect -1061 2431 -1049 2465
rect -1015 2431 -1003 2465
rect -1061 2397 -1003 2431
rect -1061 2363 -1049 2397
rect -1015 2363 -1003 2397
rect -1061 2329 -1003 2363
rect -1061 2295 -1049 2329
rect -1015 2295 -1003 2329
rect -1061 2261 -1003 2295
rect -1061 2227 -1049 2261
rect -1015 2227 -1003 2261
rect -1061 2193 -1003 2227
rect -1061 2159 -1049 2193
rect -1015 2159 -1003 2193
rect -1061 2125 -1003 2159
rect -1061 2091 -1049 2125
rect -1015 2091 -1003 2125
rect -1061 2057 -1003 2091
rect -1061 2023 -1049 2057
rect -1015 2023 -1003 2057
rect -1061 1989 -1003 2023
rect -1061 1955 -1049 1989
rect -1015 1955 -1003 1989
rect -1061 1921 -1003 1955
rect -1061 1887 -1049 1921
rect -1015 1887 -1003 1921
rect -1061 1853 -1003 1887
rect -1061 1819 -1049 1853
rect -1015 1819 -1003 1853
rect -1061 1785 -1003 1819
rect -1061 1751 -1049 1785
rect -1015 1751 -1003 1785
rect -1061 1717 -1003 1751
rect -1061 1683 -1049 1717
rect -1015 1683 -1003 1717
rect -1061 1649 -1003 1683
rect -1061 1615 -1049 1649
rect -1015 1615 -1003 1649
rect -1061 1581 -1003 1615
rect -1061 1547 -1049 1581
rect -1015 1547 -1003 1581
rect -1061 1513 -1003 1547
rect -1061 1479 -1049 1513
rect -1015 1479 -1003 1513
rect -1061 1445 -1003 1479
rect -1061 1411 -1049 1445
rect -1015 1411 -1003 1445
rect -1061 1377 -1003 1411
rect -1061 1343 -1049 1377
rect -1015 1343 -1003 1377
rect -1061 1309 -1003 1343
rect -1061 1275 -1049 1309
rect -1015 1275 -1003 1309
rect -1061 1241 -1003 1275
rect -1061 1207 -1049 1241
rect -1015 1207 -1003 1241
rect -1061 1173 -1003 1207
rect -1061 1139 -1049 1173
rect -1015 1139 -1003 1173
rect -1061 1105 -1003 1139
rect -1061 1071 -1049 1105
rect -1015 1071 -1003 1105
rect -1061 1037 -1003 1071
rect -1061 1003 -1049 1037
rect -1015 1003 -1003 1037
rect -1061 969 -1003 1003
rect -1061 935 -1049 969
rect -1015 935 -1003 969
rect -1061 901 -1003 935
rect -1061 867 -1049 901
rect -1015 867 -1003 901
rect -1061 833 -1003 867
rect -1061 799 -1049 833
rect -1015 799 -1003 833
rect -1061 765 -1003 799
rect -1061 731 -1049 765
rect -1015 731 -1003 765
rect -1061 697 -1003 731
rect -1061 663 -1049 697
rect -1015 663 -1003 697
rect -1061 629 -1003 663
rect -1061 595 -1049 629
rect -1015 595 -1003 629
rect -1061 561 -1003 595
rect -1061 527 -1049 561
rect -1015 527 -1003 561
rect -1061 493 -1003 527
rect -1061 459 -1049 493
rect -1015 459 -1003 493
rect -1061 425 -1003 459
rect -1061 391 -1049 425
rect -1015 391 -1003 425
rect -1061 357 -1003 391
rect -1061 323 -1049 357
rect -1015 323 -1003 357
rect -1061 289 -1003 323
rect -1061 255 -1049 289
rect -1015 255 -1003 289
rect -1061 221 -1003 255
rect -1061 187 -1049 221
rect -1015 187 -1003 221
rect -1061 153 -1003 187
rect -1061 119 -1049 153
rect -1015 119 -1003 153
rect -1061 85 -1003 119
rect -1061 51 -1049 85
rect -1015 51 -1003 85
rect -1061 17 -1003 51
rect -1061 -17 -1049 17
rect -1015 -17 -1003 17
rect -1061 -51 -1003 -17
rect -1061 -85 -1049 -51
rect -1015 -85 -1003 -51
rect -1061 -119 -1003 -85
rect -1061 -153 -1049 -119
rect -1015 -153 -1003 -119
rect -1061 -187 -1003 -153
rect -1061 -221 -1049 -187
rect -1015 -221 -1003 -187
rect -1061 -255 -1003 -221
rect -1061 -289 -1049 -255
rect -1015 -289 -1003 -255
rect -1061 -323 -1003 -289
rect -1061 -357 -1049 -323
rect -1015 -357 -1003 -323
rect -1061 -391 -1003 -357
rect -1061 -425 -1049 -391
rect -1015 -425 -1003 -391
rect -1061 -459 -1003 -425
rect -1061 -493 -1049 -459
rect -1015 -493 -1003 -459
rect -1061 -527 -1003 -493
rect -1061 -561 -1049 -527
rect -1015 -561 -1003 -527
rect -1061 -595 -1003 -561
rect -1061 -629 -1049 -595
rect -1015 -629 -1003 -595
rect -1061 -663 -1003 -629
rect -1061 -697 -1049 -663
rect -1015 -697 -1003 -663
rect -1061 -731 -1003 -697
rect -1061 -765 -1049 -731
rect -1015 -765 -1003 -731
rect -1061 -799 -1003 -765
rect -1061 -833 -1049 -799
rect -1015 -833 -1003 -799
rect -1061 -867 -1003 -833
rect -1061 -901 -1049 -867
rect -1015 -901 -1003 -867
rect -1061 -935 -1003 -901
rect -1061 -969 -1049 -935
rect -1015 -969 -1003 -935
rect -1061 -1003 -1003 -969
rect -1061 -1037 -1049 -1003
rect -1015 -1037 -1003 -1003
rect -1061 -1071 -1003 -1037
rect -1061 -1105 -1049 -1071
rect -1015 -1105 -1003 -1071
rect -1061 -1139 -1003 -1105
rect -1061 -1173 -1049 -1139
rect -1015 -1173 -1003 -1139
rect -1061 -1207 -1003 -1173
rect -1061 -1241 -1049 -1207
rect -1015 -1241 -1003 -1207
rect -1061 -1275 -1003 -1241
rect -1061 -1309 -1049 -1275
rect -1015 -1309 -1003 -1275
rect -1061 -1343 -1003 -1309
rect -1061 -1377 -1049 -1343
rect -1015 -1377 -1003 -1343
rect -1061 -1411 -1003 -1377
rect -1061 -1445 -1049 -1411
rect -1015 -1445 -1003 -1411
rect -1061 -1479 -1003 -1445
rect -1061 -1513 -1049 -1479
rect -1015 -1513 -1003 -1479
rect -1061 -1547 -1003 -1513
rect -1061 -1581 -1049 -1547
rect -1015 -1581 -1003 -1547
rect -1061 -1615 -1003 -1581
rect -1061 -1649 -1049 -1615
rect -1015 -1649 -1003 -1615
rect -1061 -1683 -1003 -1649
rect -1061 -1717 -1049 -1683
rect -1015 -1717 -1003 -1683
rect -1061 -1751 -1003 -1717
rect -1061 -1785 -1049 -1751
rect -1015 -1785 -1003 -1751
rect -1061 -1819 -1003 -1785
rect -1061 -1853 -1049 -1819
rect -1015 -1853 -1003 -1819
rect -1061 -1887 -1003 -1853
rect -1061 -1921 -1049 -1887
rect -1015 -1921 -1003 -1887
rect -1061 -1955 -1003 -1921
rect -1061 -1989 -1049 -1955
rect -1015 -1989 -1003 -1955
rect -1061 -2023 -1003 -1989
rect -1061 -2057 -1049 -2023
rect -1015 -2057 -1003 -2023
rect -1061 -2091 -1003 -2057
rect -1061 -2125 -1049 -2091
rect -1015 -2125 -1003 -2091
rect -1061 -2159 -1003 -2125
rect -1061 -2193 -1049 -2159
rect -1015 -2193 -1003 -2159
rect -1061 -2227 -1003 -2193
rect -1061 -2261 -1049 -2227
rect -1015 -2261 -1003 -2227
rect -1061 -2295 -1003 -2261
rect -1061 -2329 -1049 -2295
rect -1015 -2329 -1003 -2295
rect -1061 -2363 -1003 -2329
rect -1061 -2397 -1049 -2363
rect -1015 -2397 -1003 -2363
rect -1061 -2431 -1003 -2397
rect -1061 -2465 -1049 -2431
rect -1015 -2465 -1003 -2431
rect -1061 -2500 -1003 -2465
rect -803 2465 -745 2500
rect -803 2431 -791 2465
rect -757 2431 -745 2465
rect -803 2397 -745 2431
rect -803 2363 -791 2397
rect -757 2363 -745 2397
rect -803 2329 -745 2363
rect -803 2295 -791 2329
rect -757 2295 -745 2329
rect -803 2261 -745 2295
rect -803 2227 -791 2261
rect -757 2227 -745 2261
rect -803 2193 -745 2227
rect -803 2159 -791 2193
rect -757 2159 -745 2193
rect -803 2125 -745 2159
rect -803 2091 -791 2125
rect -757 2091 -745 2125
rect -803 2057 -745 2091
rect -803 2023 -791 2057
rect -757 2023 -745 2057
rect -803 1989 -745 2023
rect -803 1955 -791 1989
rect -757 1955 -745 1989
rect -803 1921 -745 1955
rect -803 1887 -791 1921
rect -757 1887 -745 1921
rect -803 1853 -745 1887
rect -803 1819 -791 1853
rect -757 1819 -745 1853
rect -803 1785 -745 1819
rect -803 1751 -791 1785
rect -757 1751 -745 1785
rect -803 1717 -745 1751
rect -803 1683 -791 1717
rect -757 1683 -745 1717
rect -803 1649 -745 1683
rect -803 1615 -791 1649
rect -757 1615 -745 1649
rect -803 1581 -745 1615
rect -803 1547 -791 1581
rect -757 1547 -745 1581
rect -803 1513 -745 1547
rect -803 1479 -791 1513
rect -757 1479 -745 1513
rect -803 1445 -745 1479
rect -803 1411 -791 1445
rect -757 1411 -745 1445
rect -803 1377 -745 1411
rect -803 1343 -791 1377
rect -757 1343 -745 1377
rect -803 1309 -745 1343
rect -803 1275 -791 1309
rect -757 1275 -745 1309
rect -803 1241 -745 1275
rect -803 1207 -791 1241
rect -757 1207 -745 1241
rect -803 1173 -745 1207
rect -803 1139 -791 1173
rect -757 1139 -745 1173
rect -803 1105 -745 1139
rect -803 1071 -791 1105
rect -757 1071 -745 1105
rect -803 1037 -745 1071
rect -803 1003 -791 1037
rect -757 1003 -745 1037
rect -803 969 -745 1003
rect -803 935 -791 969
rect -757 935 -745 969
rect -803 901 -745 935
rect -803 867 -791 901
rect -757 867 -745 901
rect -803 833 -745 867
rect -803 799 -791 833
rect -757 799 -745 833
rect -803 765 -745 799
rect -803 731 -791 765
rect -757 731 -745 765
rect -803 697 -745 731
rect -803 663 -791 697
rect -757 663 -745 697
rect -803 629 -745 663
rect -803 595 -791 629
rect -757 595 -745 629
rect -803 561 -745 595
rect -803 527 -791 561
rect -757 527 -745 561
rect -803 493 -745 527
rect -803 459 -791 493
rect -757 459 -745 493
rect -803 425 -745 459
rect -803 391 -791 425
rect -757 391 -745 425
rect -803 357 -745 391
rect -803 323 -791 357
rect -757 323 -745 357
rect -803 289 -745 323
rect -803 255 -791 289
rect -757 255 -745 289
rect -803 221 -745 255
rect -803 187 -791 221
rect -757 187 -745 221
rect -803 153 -745 187
rect -803 119 -791 153
rect -757 119 -745 153
rect -803 85 -745 119
rect -803 51 -791 85
rect -757 51 -745 85
rect -803 17 -745 51
rect -803 -17 -791 17
rect -757 -17 -745 17
rect -803 -51 -745 -17
rect -803 -85 -791 -51
rect -757 -85 -745 -51
rect -803 -119 -745 -85
rect -803 -153 -791 -119
rect -757 -153 -745 -119
rect -803 -187 -745 -153
rect -803 -221 -791 -187
rect -757 -221 -745 -187
rect -803 -255 -745 -221
rect -803 -289 -791 -255
rect -757 -289 -745 -255
rect -803 -323 -745 -289
rect -803 -357 -791 -323
rect -757 -357 -745 -323
rect -803 -391 -745 -357
rect -803 -425 -791 -391
rect -757 -425 -745 -391
rect -803 -459 -745 -425
rect -803 -493 -791 -459
rect -757 -493 -745 -459
rect -803 -527 -745 -493
rect -803 -561 -791 -527
rect -757 -561 -745 -527
rect -803 -595 -745 -561
rect -803 -629 -791 -595
rect -757 -629 -745 -595
rect -803 -663 -745 -629
rect -803 -697 -791 -663
rect -757 -697 -745 -663
rect -803 -731 -745 -697
rect -803 -765 -791 -731
rect -757 -765 -745 -731
rect -803 -799 -745 -765
rect -803 -833 -791 -799
rect -757 -833 -745 -799
rect -803 -867 -745 -833
rect -803 -901 -791 -867
rect -757 -901 -745 -867
rect -803 -935 -745 -901
rect -803 -969 -791 -935
rect -757 -969 -745 -935
rect -803 -1003 -745 -969
rect -803 -1037 -791 -1003
rect -757 -1037 -745 -1003
rect -803 -1071 -745 -1037
rect -803 -1105 -791 -1071
rect -757 -1105 -745 -1071
rect -803 -1139 -745 -1105
rect -803 -1173 -791 -1139
rect -757 -1173 -745 -1139
rect -803 -1207 -745 -1173
rect -803 -1241 -791 -1207
rect -757 -1241 -745 -1207
rect -803 -1275 -745 -1241
rect -803 -1309 -791 -1275
rect -757 -1309 -745 -1275
rect -803 -1343 -745 -1309
rect -803 -1377 -791 -1343
rect -757 -1377 -745 -1343
rect -803 -1411 -745 -1377
rect -803 -1445 -791 -1411
rect -757 -1445 -745 -1411
rect -803 -1479 -745 -1445
rect -803 -1513 -791 -1479
rect -757 -1513 -745 -1479
rect -803 -1547 -745 -1513
rect -803 -1581 -791 -1547
rect -757 -1581 -745 -1547
rect -803 -1615 -745 -1581
rect -803 -1649 -791 -1615
rect -757 -1649 -745 -1615
rect -803 -1683 -745 -1649
rect -803 -1717 -791 -1683
rect -757 -1717 -745 -1683
rect -803 -1751 -745 -1717
rect -803 -1785 -791 -1751
rect -757 -1785 -745 -1751
rect -803 -1819 -745 -1785
rect -803 -1853 -791 -1819
rect -757 -1853 -745 -1819
rect -803 -1887 -745 -1853
rect -803 -1921 -791 -1887
rect -757 -1921 -745 -1887
rect -803 -1955 -745 -1921
rect -803 -1989 -791 -1955
rect -757 -1989 -745 -1955
rect -803 -2023 -745 -1989
rect -803 -2057 -791 -2023
rect -757 -2057 -745 -2023
rect -803 -2091 -745 -2057
rect -803 -2125 -791 -2091
rect -757 -2125 -745 -2091
rect -803 -2159 -745 -2125
rect -803 -2193 -791 -2159
rect -757 -2193 -745 -2159
rect -803 -2227 -745 -2193
rect -803 -2261 -791 -2227
rect -757 -2261 -745 -2227
rect -803 -2295 -745 -2261
rect -803 -2329 -791 -2295
rect -757 -2329 -745 -2295
rect -803 -2363 -745 -2329
rect -803 -2397 -791 -2363
rect -757 -2397 -745 -2363
rect -803 -2431 -745 -2397
rect -803 -2465 -791 -2431
rect -757 -2465 -745 -2431
rect -803 -2500 -745 -2465
rect -545 2465 -487 2500
rect -545 2431 -533 2465
rect -499 2431 -487 2465
rect -545 2397 -487 2431
rect -545 2363 -533 2397
rect -499 2363 -487 2397
rect -545 2329 -487 2363
rect -545 2295 -533 2329
rect -499 2295 -487 2329
rect -545 2261 -487 2295
rect -545 2227 -533 2261
rect -499 2227 -487 2261
rect -545 2193 -487 2227
rect -545 2159 -533 2193
rect -499 2159 -487 2193
rect -545 2125 -487 2159
rect -545 2091 -533 2125
rect -499 2091 -487 2125
rect -545 2057 -487 2091
rect -545 2023 -533 2057
rect -499 2023 -487 2057
rect -545 1989 -487 2023
rect -545 1955 -533 1989
rect -499 1955 -487 1989
rect -545 1921 -487 1955
rect -545 1887 -533 1921
rect -499 1887 -487 1921
rect -545 1853 -487 1887
rect -545 1819 -533 1853
rect -499 1819 -487 1853
rect -545 1785 -487 1819
rect -545 1751 -533 1785
rect -499 1751 -487 1785
rect -545 1717 -487 1751
rect -545 1683 -533 1717
rect -499 1683 -487 1717
rect -545 1649 -487 1683
rect -545 1615 -533 1649
rect -499 1615 -487 1649
rect -545 1581 -487 1615
rect -545 1547 -533 1581
rect -499 1547 -487 1581
rect -545 1513 -487 1547
rect -545 1479 -533 1513
rect -499 1479 -487 1513
rect -545 1445 -487 1479
rect -545 1411 -533 1445
rect -499 1411 -487 1445
rect -545 1377 -487 1411
rect -545 1343 -533 1377
rect -499 1343 -487 1377
rect -545 1309 -487 1343
rect -545 1275 -533 1309
rect -499 1275 -487 1309
rect -545 1241 -487 1275
rect -545 1207 -533 1241
rect -499 1207 -487 1241
rect -545 1173 -487 1207
rect -545 1139 -533 1173
rect -499 1139 -487 1173
rect -545 1105 -487 1139
rect -545 1071 -533 1105
rect -499 1071 -487 1105
rect -545 1037 -487 1071
rect -545 1003 -533 1037
rect -499 1003 -487 1037
rect -545 969 -487 1003
rect -545 935 -533 969
rect -499 935 -487 969
rect -545 901 -487 935
rect -545 867 -533 901
rect -499 867 -487 901
rect -545 833 -487 867
rect -545 799 -533 833
rect -499 799 -487 833
rect -545 765 -487 799
rect -545 731 -533 765
rect -499 731 -487 765
rect -545 697 -487 731
rect -545 663 -533 697
rect -499 663 -487 697
rect -545 629 -487 663
rect -545 595 -533 629
rect -499 595 -487 629
rect -545 561 -487 595
rect -545 527 -533 561
rect -499 527 -487 561
rect -545 493 -487 527
rect -545 459 -533 493
rect -499 459 -487 493
rect -545 425 -487 459
rect -545 391 -533 425
rect -499 391 -487 425
rect -545 357 -487 391
rect -545 323 -533 357
rect -499 323 -487 357
rect -545 289 -487 323
rect -545 255 -533 289
rect -499 255 -487 289
rect -545 221 -487 255
rect -545 187 -533 221
rect -499 187 -487 221
rect -545 153 -487 187
rect -545 119 -533 153
rect -499 119 -487 153
rect -545 85 -487 119
rect -545 51 -533 85
rect -499 51 -487 85
rect -545 17 -487 51
rect -545 -17 -533 17
rect -499 -17 -487 17
rect -545 -51 -487 -17
rect -545 -85 -533 -51
rect -499 -85 -487 -51
rect -545 -119 -487 -85
rect -545 -153 -533 -119
rect -499 -153 -487 -119
rect -545 -187 -487 -153
rect -545 -221 -533 -187
rect -499 -221 -487 -187
rect -545 -255 -487 -221
rect -545 -289 -533 -255
rect -499 -289 -487 -255
rect -545 -323 -487 -289
rect -545 -357 -533 -323
rect -499 -357 -487 -323
rect -545 -391 -487 -357
rect -545 -425 -533 -391
rect -499 -425 -487 -391
rect -545 -459 -487 -425
rect -545 -493 -533 -459
rect -499 -493 -487 -459
rect -545 -527 -487 -493
rect -545 -561 -533 -527
rect -499 -561 -487 -527
rect -545 -595 -487 -561
rect -545 -629 -533 -595
rect -499 -629 -487 -595
rect -545 -663 -487 -629
rect -545 -697 -533 -663
rect -499 -697 -487 -663
rect -545 -731 -487 -697
rect -545 -765 -533 -731
rect -499 -765 -487 -731
rect -545 -799 -487 -765
rect -545 -833 -533 -799
rect -499 -833 -487 -799
rect -545 -867 -487 -833
rect -545 -901 -533 -867
rect -499 -901 -487 -867
rect -545 -935 -487 -901
rect -545 -969 -533 -935
rect -499 -969 -487 -935
rect -545 -1003 -487 -969
rect -545 -1037 -533 -1003
rect -499 -1037 -487 -1003
rect -545 -1071 -487 -1037
rect -545 -1105 -533 -1071
rect -499 -1105 -487 -1071
rect -545 -1139 -487 -1105
rect -545 -1173 -533 -1139
rect -499 -1173 -487 -1139
rect -545 -1207 -487 -1173
rect -545 -1241 -533 -1207
rect -499 -1241 -487 -1207
rect -545 -1275 -487 -1241
rect -545 -1309 -533 -1275
rect -499 -1309 -487 -1275
rect -545 -1343 -487 -1309
rect -545 -1377 -533 -1343
rect -499 -1377 -487 -1343
rect -545 -1411 -487 -1377
rect -545 -1445 -533 -1411
rect -499 -1445 -487 -1411
rect -545 -1479 -487 -1445
rect -545 -1513 -533 -1479
rect -499 -1513 -487 -1479
rect -545 -1547 -487 -1513
rect -545 -1581 -533 -1547
rect -499 -1581 -487 -1547
rect -545 -1615 -487 -1581
rect -545 -1649 -533 -1615
rect -499 -1649 -487 -1615
rect -545 -1683 -487 -1649
rect -545 -1717 -533 -1683
rect -499 -1717 -487 -1683
rect -545 -1751 -487 -1717
rect -545 -1785 -533 -1751
rect -499 -1785 -487 -1751
rect -545 -1819 -487 -1785
rect -545 -1853 -533 -1819
rect -499 -1853 -487 -1819
rect -545 -1887 -487 -1853
rect -545 -1921 -533 -1887
rect -499 -1921 -487 -1887
rect -545 -1955 -487 -1921
rect -545 -1989 -533 -1955
rect -499 -1989 -487 -1955
rect -545 -2023 -487 -1989
rect -545 -2057 -533 -2023
rect -499 -2057 -487 -2023
rect -545 -2091 -487 -2057
rect -545 -2125 -533 -2091
rect -499 -2125 -487 -2091
rect -545 -2159 -487 -2125
rect -545 -2193 -533 -2159
rect -499 -2193 -487 -2159
rect -545 -2227 -487 -2193
rect -545 -2261 -533 -2227
rect -499 -2261 -487 -2227
rect -545 -2295 -487 -2261
rect -545 -2329 -533 -2295
rect -499 -2329 -487 -2295
rect -545 -2363 -487 -2329
rect -545 -2397 -533 -2363
rect -499 -2397 -487 -2363
rect -545 -2431 -487 -2397
rect -545 -2465 -533 -2431
rect -499 -2465 -487 -2431
rect -545 -2500 -487 -2465
rect -287 2465 -229 2500
rect -287 2431 -275 2465
rect -241 2431 -229 2465
rect -287 2397 -229 2431
rect -287 2363 -275 2397
rect -241 2363 -229 2397
rect -287 2329 -229 2363
rect -287 2295 -275 2329
rect -241 2295 -229 2329
rect -287 2261 -229 2295
rect -287 2227 -275 2261
rect -241 2227 -229 2261
rect -287 2193 -229 2227
rect -287 2159 -275 2193
rect -241 2159 -229 2193
rect -287 2125 -229 2159
rect -287 2091 -275 2125
rect -241 2091 -229 2125
rect -287 2057 -229 2091
rect -287 2023 -275 2057
rect -241 2023 -229 2057
rect -287 1989 -229 2023
rect -287 1955 -275 1989
rect -241 1955 -229 1989
rect -287 1921 -229 1955
rect -287 1887 -275 1921
rect -241 1887 -229 1921
rect -287 1853 -229 1887
rect -287 1819 -275 1853
rect -241 1819 -229 1853
rect -287 1785 -229 1819
rect -287 1751 -275 1785
rect -241 1751 -229 1785
rect -287 1717 -229 1751
rect -287 1683 -275 1717
rect -241 1683 -229 1717
rect -287 1649 -229 1683
rect -287 1615 -275 1649
rect -241 1615 -229 1649
rect -287 1581 -229 1615
rect -287 1547 -275 1581
rect -241 1547 -229 1581
rect -287 1513 -229 1547
rect -287 1479 -275 1513
rect -241 1479 -229 1513
rect -287 1445 -229 1479
rect -287 1411 -275 1445
rect -241 1411 -229 1445
rect -287 1377 -229 1411
rect -287 1343 -275 1377
rect -241 1343 -229 1377
rect -287 1309 -229 1343
rect -287 1275 -275 1309
rect -241 1275 -229 1309
rect -287 1241 -229 1275
rect -287 1207 -275 1241
rect -241 1207 -229 1241
rect -287 1173 -229 1207
rect -287 1139 -275 1173
rect -241 1139 -229 1173
rect -287 1105 -229 1139
rect -287 1071 -275 1105
rect -241 1071 -229 1105
rect -287 1037 -229 1071
rect -287 1003 -275 1037
rect -241 1003 -229 1037
rect -287 969 -229 1003
rect -287 935 -275 969
rect -241 935 -229 969
rect -287 901 -229 935
rect -287 867 -275 901
rect -241 867 -229 901
rect -287 833 -229 867
rect -287 799 -275 833
rect -241 799 -229 833
rect -287 765 -229 799
rect -287 731 -275 765
rect -241 731 -229 765
rect -287 697 -229 731
rect -287 663 -275 697
rect -241 663 -229 697
rect -287 629 -229 663
rect -287 595 -275 629
rect -241 595 -229 629
rect -287 561 -229 595
rect -287 527 -275 561
rect -241 527 -229 561
rect -287 493 -229 527
rect -287 459 -275 493
rect -241 459 -229 493
rect -287 425 -229 459
rect -287 391 -275 425
rect -241 391 -229 425
rect -287 357 -229 391
rect -287 323 -275 357
rect -241 323 -229 357
rect -287 289 -229 323
rect -287 255 -275 289
rect -241 255 -229 289
rect -287 221 -229 255
rect -287 187 -275 221
rect -241 187 -229 221
rect -287 153 -229 187
rect -287 119 -275 153
rect -241 119 -229 153
rect -287 85 -229 119
rect -287 51 -275 85
rect -241 51 -229 85
rect -287 17 -229 51
rect -287 -17 -275 17
rect -241 -17 -229 17
rect -287 -51 -229 -17
rect -287 -85 -275 -51
rect -241 -85 -229 -51
rect -287 -119 -229 -85
rect -287 -153 -275 -119
rect -241 -153 -229 -119
rect -287 -187 -229 -153
rect -287 -221 -275 -187
rect -241 -221 -229 -187
rect -287 -255 -229 -221
rect -287 -289 -275 -255
rect -241 -289 -229 -255
rect -287 -323 -229 -289
rect -287 -357 -275 -323
rect -241 -357 -229 -323
rect -287 -391 -229 -357
rect -287 -425 -275 -391
rect -241 -425 -229 -391
rect -287 -459 -229 -425
rect -287 -493 -275 -459
rect -241 -493 -229 -459
rect -287 -527 -229 -493
rect -287 -561 -275 -527
rect -241 -561 -229 -527
rect -287 -595 -229 -561
rect -287 -629 -275 -595
rect -241 -629 -229 -595
rect -287 -663 -229 -629
rect -287 -697 -275 -663
rect -241 -697 -229 -663
rect -287 -731 -229 -697
rect -287 -765 -275 -731
rect -241 -765 -229 -731
rect -287 -799 -229 -765
rect -287 -833 -275 -799
rect -241 -833 -229 -799
rect -287 -867 -229 -833
rect -287 -901 -275 -867
rect -241 -901 -229 -867
rect -287 -935 -229 -901
rect -287 -969 -275 -935
rect -241 -969 -229 -935
rect -287 -1003 -229 -969
rect -287 -1037 -275 -1003
rect -241 -1037 -229 -1003
rect -287 -1071 -229 -1037
rect -287 -1105 -275 -1071
rect -241 -1105 -229 -1071
rect -287 -1139 -229 -1105
rect -287 -1173 -275 -1139
rect -241 -1173 -229 -1139
rect -287 -1207 -229 -1173
rect -287 -1241 -275 -1207
rect -241 -1241 -229 -1207
rect -287 -1275 -229 -1241
rect -287 -1309 -275 -1275
rect -241 -1309 -229 -1275
rect -287 -1343 -229 -1309
rect -287 -1377 -275 -1343
rect -241 -1377 -229 -1343
rect -287 -1411 -229 -1377
rect -287 -1445 -275 -1411
rect -241 -1445 -229 -1411
rect -287 -1479 -229 -1445
rect -287 -1513 -275 -1479
rect -241 -1513 -229 -1479
rect -287 -1547 -229 -1513
rect -287 -1581 -275 -1547
rect -241 -1581 -229 -1547
rect -287 -1615 -229 -1581
rect -287 -1649 -275 -1615
rect -241 -1649 -229 -1615
rect -287 -1683 -229 -1649
rect -287 -1717 -275 -1683
rect -241 -1717 -229 -1683
rect -287 -1751 -229 -1717
rect -287 -1785 -275 -1751
rect -241 -1785 -229 -1751
rect -287 -1819 -229 -1785
rect -287 -1853 -275 -1819
rect -241 -1853 -229 -1819
rect -287 -1887 -229 -1853
rect -287 -1921 -275 -1887
rect -241 -1921 -229 -1887
rect -287 -1955 -229 -1921
rect -287 -1989 -275 -1955
rect -241 -1989 -229 -1955
rect -287 -2023 -229 -1989
rect -287 -2057 -275 -2023
rect -241 -2057 -229 -2023
rect -287 -2091 -229 -2057
rect -287 -2125 -275 -2091
rect -241 -2125 -229 -2091
rect -287 -2159 -229 -2125
rect -287 -2193 -275 -2159
rect -241 -2193 -229 -2159
rect -287 -2227 -229 -2193
rect -287 -2261 -275 -2227
rect -241 -2261 -229 -2227
rect -287 -2295 -229 -2261
rect -287 -2329 -275 -2295
rect -241 -2329 -229 -2295
rect -287 -2363 -229 -2329
rect -287 -2397 -275 -2363
rect -241 -2397 -229 -2363
rect -287 -2431 -229 -2397
rect -287 -2465 -275 -2431
rect -241 -2465 -229 -2431
rect -287 -2500 -229 -2465
rect -29 2465 29 2500
rect -29 2431 -17 2465
rect 17 2431 29 2465
rect -29 2397 29 2431
rect -29 2363 -17 2397
rect 17 2363 29 2397
rect -29 2329 29 2363
rect -29 2295 -17 2329
rect 17 2295 29 2329
rect -29 2261 29 2295
rect -29 2227 -17 2261
rect 17 2227 29 2261
rect -29 2193 29 2227
rect -29 2159 -17 2193
rect 17 2159 29 2193
rect -29 2125 29 2159
rect -29 2091 -17 2125
rect 17 2091 29 2125
rect -29 2057 29 2091
rect -29 2023 -17 2057
rect 17 2023 29 2057
rect -29 1989 29 2023
rect -29 1955 -17 1989
rect 17 1955 29 1989
rect -29 1921 29 1955
rect -29 1887 -17 1921
rect 17 1887 29 1921
rect -29 1853 29 1887
rect -29 1819 -17 1853
rect 17 1819 29 1853
rect -29 1785 29 1819
rect -29 1751 -17 1785
rect 17 1751 29 1785
rect -29 1717 29 1751
rect -29 1683 -17 1717
rect 17 1683 29 1717
rect -29 1649 29 1683
rect -29 1615 -17 1649
rect 17 1615 29 1649
rect -29 1581 29 1615
rect -29 1547 -17 1581
rect 17 1547 29 1581
rect -29 1513 29 1547
rect -29 1479 -17 1513
rect 17 1479 29 1513
rect -29 1445 29 1479
rect -29 1411 -17 1445
rect 17 1411 29 1445
rect -29 1377 29 1411
rect -29 1343 -17 1377
rect 17 1343 29 1377
rect -29 1309 29 1343
rect -29 1275 -17 1309
rect 17 1275 29 1309
rect -29 1241 29 1275
rect -29 1207 -17 1241
rect 17 1207 29 1241
rect -29 1173 29 1207
rect -29 1139 -17 1173
rect 17 1139 29 1173
rect -29 1105 29 1139
rect -29 1071 -17 1105
rect 17 1071 29 1105
rect -29 1037 29 1071
rect -29 1003 -17 1037
rect 17 1003 29 1037
rect -29 969 29 1003
rect -29 935 -17 969
rect 17 935 29 969
rect -29 901 29 935
rect -29 867 -17 901
rect 17 867 29 901
rect -29 833 29 867
rect -29 799 -17 833
rect 17 799 29 833
rect -29 765 29 799
rect -29 731 -17 765
rect 17 731 29 765
rect -29 697 29 731
rect -29 663 -17 697
rect 17 663 29 697
rect -29 629 29 663
rect -29 595 -17 629
rect 17 595 29 629
rect -29 561 29 595
rect -29 527 -17 561
rect 17 527 29 561
rect -29 493 29 527
rect -29 459 -17 493
rect 17 459 29 493
rect -29 425 29 459
rect -29 391 -17 425
rect 17 391 29 425
rect -29 357 29 391
rect -29 323 -17 357
rect 17 323 29 357
rect -29 289 29 323
rect -29 255 -17 289
rect 17 255 29 289
rect -29 221 29 255
rect -29 187 -17 221
rect 17 187 29 221
rect -29 153 29 187
rect -29 119 -17 153
rect 17 119 29 153
rect -29 85 29 119
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -119 29 -85
rect -29 -153 -17 -119
rect 17 -153 29 -119
rect -29 -187 29 -153
rect -29 -221 -17 -187
rect 17 -221 29 -187
rect -29 -255 29 -221
rect -29 -289 -17 -255
rect 17 -289 29 -255
rect -29 -323 29 -289
rect -29 -357 -17 -323
rect 17 -357 29 -323
rect -29 -391 29 -357
rect -29 -425 -17 -391
rect 17 -425 29 -391
rect -29 -459 29 -425
rect -29 -493 -17 -459
rect 17 -493 29 -459
rect -29 -527 29 -493
rect -29 -561 -17 -527
rect 17 -561 29 -527
rect -29 -595 29 -561
rect -29 -629 -17 -595
rect 17 -629 29 -595
rect -29 -663 29 -629
rect -29 -697 -17 -663
rect 17 -697 29 -663
rect -29 -731 29 -697
rect -29 -765 -17 -731
rect 17 -765 29 -731
rect -29 -799 29 -765
rect -29 -833 -17 -799
rect 17 -833 29 -799
rect -29 -867 29 -833
rect -29 -901 -17 -867
rect 17 -901 29 -867
rect -29 -935 29 -901
rect -29 -969 -17 -935
rect 17 -969 29 -935
rect -29 -1003 29 -969
rect -29 -1037 -17 -1003
rect 17 -1037 29 -1003
rect -29 -1071 29 -1037
rect -29 -1105 -17 -1071
rect 17 -1105 29 -1071
rect -29 -1139 29 -1105
rect -29 -1173 -17 -1139
rect 17 -1173 29 -1139
rect -29 -1207 29 -1173
rect -29 -1241 -17 -1207
rect 17 -1241 29 -1207
rect -29 -1275 29 -1241
rect -29 -1309 -17 -1275
rect 17 -1309 29 -1275
rect -29 -1343 29 -1309
rect -29 -1377 -17 -1343
rect 17 -1377 29 -1343
rect -29 -1411 29 -1377
rect -29 -1445 -17 -1411
rect 17 -1445 29 -1411
rect -29 -1479 29 -1445
rect -29 -1513 -17 -1479
rect 17 -1513 29 -1479
rect -29 -1547 29 -1513
rect -29 -1581 -17 -1547
rect 17 -1581 29 -1547
rect -29 -1615 29 -1581
rect -29 -1649 -17 -1615
rect 17 -1649 29 -1615
rect -29 -1683 29 -1649
rect -29 -1717 -17 -1683
rect 17 -1717 29 -1683
rect -29 -1751 29 -1717
rect -29 -1785 -17 -1751
rect 17 -1785 29 -1751
rect -29 -1819 29 -1785
rect -29 -1853 -17 -1819
rect 17 -1853 29 -1819
rect -29 -1887 29 -1853
rect -29 -1921 -17 -1887
rect 17 -1921 29 -1887
rect -29 -1955 29 -1921
rect -29 -1989 -17 -1955
rect 17 -1989 29 -1955
rect -29 -2023 29 -1989
rect -29 -2057 -17 -2023
rect 17 -2057 29 -2023
rect -29 -2091 29 -2057
rect -29 -2125 -17 -2091
rect 17 -2125 29 -2091
rect -29 -2159 29 -2125
rect -29 -2193 -17 -2159
rect 17 -2193 29 -2159
rect -29 -2227 29 -2193
rect -29 -2261 -17 -2227
rect 17 -2261 29 -2227
rect -29 -2295 29 -2261
rect -29 -2329 -17 -2295
rect 17 -2329 29 -2295
rect -29 -2363 29 -2329
rect -29 -2397 -17 -2363
rect 17 -2397 29 -2363
rect -29 -2431 29 -2397
rect -29 -2465 -17 -2431
rect 17 -2465 29 -2431
rect -29 -2500 29 -2465
rect 229 2465 287 2500
rect 229 2431 241 2465
rect 275 2431 287 2465
rect 229 2397 287 2431
rect 229 2363 241 2397
rect 275 2363 287 2397
rect 229 2329 287 2363
rect 229 2295 241 2329
rect 275 2295 287 2329
rect 229 2261 287 2295
rect 229 2227 241 2261
rect 275 2227 287 2261
rect 229 2193 287 2227
rect 229 2159 241 2193
rect 275 2159 287 2193
rect 229 2125 287 2159
rect 229 2091 241 2125
rect 275 2091 287 2125
rect 229 2057 287 2091
rect 229 2023 241 2057
rect 275 2023 287 2057
rect 229 1989 287 2023
rect 229 1955 241 1989
rect 275 1955 287 1989
rect 229 1921 287 1955
rect 229 1887 241 1921
rect 275 1887 287 1921
rect 229 1853 287 1887
rect 229 1819 241 1853
rect 275 1819 287 1853
rect 229 1785 287 1819
rect 229 1751 241 1785
rect 275 1751 287 1785
rect 229 1717 287 1751
rect 229 1683 241 1717
rect 275 1683 287 1717
rect 229 1649 287 1683
rect 229 1615 241 1649
rect 275 1615 287 1649
rect 229 1581 287 1615
rect 229 1547 241 1581
rect 275 1547 287 1581
rect 229 1513 287 1547
rect 229 1479 241 1513
rect 275 1479 287 1513
rect 229 1445 287 1479
rect 229 1411 241 1445
rect 275 1411 287 1445
rect 229 1377 287 1411
rect 229 1343 241 1377
rect 275 1343 287 1377
rect 229 1309 287 1343
rect 229 1275 241 1309
rect 275 1275 287 1309
rect 229 1241 287 1275
rect 229 1207 241 1241
rect 275 1207 287 1241
rect 229 1173 287 1207
rect 229 1139 241 1173
rect 275 1139 287 1173
rect 229 1105 287 1139
rect 229 1071 241 1105
rect 275 1071 287 1105
rect 229 1037 287 1071
rect 229 1003 241 1037
rect 275 1003 287 1037
rect 229 969 287 1003
rect 229 935 241 969
rect 275 935 287 969
rect 229 901 287 935
rect 229 867 241 901
rect 275 867 287 901
rect 229 833 287 867
rect 229 799 241 833
rect 275 799 287 833
rect 229 765 287 799
rect 229 731 241 765
rect 275 731 287 765
rect 229 697 287 731
rect 229 663 241 697
rect 275 663 287 697
rect 229 629 287 663
rect 229 595 241 629
rect 275 595 287 629
rect 229 561 287 595
rect 229 527 241 561
rect 275 527 287 561
rect 229 493 287 527
rect 229 459 241 493
rect 275 459 287 493
rect 229 425 287 459
rect 229 391 241 425
rect 275 391 287 425
rect 229 357 287 391
rect 229 323 241 357
rect 275 323 287 357
rect 229 289 287 323
rect 229 255 241 289
rect 275 255 287 289
rect 229 221 287 255
rect 229 187 241 221
rect 275 187 287 221
rect 229 153 287 187
rect 229 119 241 153
rect 275 119 287 153
rect 229 85 287 119
rect 229 51 241 85
rect 275 51 287 85
rect 229 17 287 51
rect 229 -17 241 17
rect 275 -17 287 17
rect 229 -51 287 -17
rect 229 -85 241 -51
rect 275 -85 287 -51
rect 229 -119 287 -85
rect 229 -153 241 -119
rect 275 -153 287 -119
rect 229 -187 287 -153
rect 229 -221 241 -187
rect 275 -221 287 -187
rect 229 -255 287 -221
rect 229 -289 241 -255
rect 275 -289 287 -255
rect 229 -323 287 -289
rect 229 -357 241 -323
rect 275 -357 287 -323
rect 229 -391 287 -357
rect 229 -425 241 -391
rect 275 -425 287 -391
rect 229 -459 287 -425
rect 229 -493 241 -459
rect 275 -493 287 -459
rect 229 -527 287 -493
rect 229 -561 241 -527
rect 275 -561 287 -527
rect 229 -595 287 -561
rect 229 -629 241 -595
rect 275 -629 287 -595
rect 229 -663 287 -629
rect 229 -697 241 -663
rect 275 -697 287 -663
rect 229 -731 287 -697
rect 229 -765 241 -731
rect 275 -765 287 -731
rect 229 -799 287 -765
rect 229 -833 241 -799
rect 275 -833 287 -799
rect 229 -867 287 -833
rect 229 -901 241 -867
rect 275 -901 287 -867
rect 229 -935 287 -901
rect 229 -969 241 -935
rect 275 -969 287 -935
rect 229 -1003 287 -969
rect 229 -1037 241 -1003
rect 275 -1037 287 -1003
rect 229 -1071 287 -1037
rect 229 -1105 241 -1071
rect 275 -1105 287 -1071
rect 229 -1139 287 -1105
rect 229 -1173 241 -1139
rect 275 -1173 287 -1139
rect 229 -1207 287 -1173
rect 229 -1241 241 -1207
rect 275 -1241 287 -1207
rect 229 -1275 287 -1241
rect 229 -1309 241 -1275
rect 275 -1309 287 -1275
rect 229 -1343 287 -1309
rect 229 -1377 241 -1343
rect 275 -1377 287 -1343
rect 229 -1411 287 -1377
rect 229 -1445 241 -1411
rect 275 -1445 287 -1411
rect 229 -1479 287 -1445
rect 229 -1513 241 -1479
rect 275 -1513 287 -1479
rect 229 -1547 287 -1513
rect 229 -1581 241 -1547
rect 275 -1581 287 -1547
rect 229 -1615 287 -1581
rect 229 -1649 241 -1615
rect 275 -1649 287 -1615
rect 229 -1683 287 -1649
rect 229 -1717 241 -1683
rect 275 -1717 287 -1683
rect 229 -1751 287 -1717
rect 229 -1785 241 -1751
rect 275 -1785 287 -1751
rect 229 -1819 287 -1785
rect 229 -1853 241 -1819
rect 275 -1853 287 -1819
rect 229 -1887 287 -1853
rect 229 -1921 241 -1887
rect 275 -1921 287 -1887
rect 229 -1955 287 -1921
rect 229 -1989 241 -1955
rect 275 -1989 287 -1955
rect 229 -2023 287 -1989
rect 229 -2057 241 -2023
rect 275 -2057 287 -2023
rect 229 -2091 287 -2057
rect 229 -2125 241 -2091
rect 275 -2125 287 -2091
rect 229 -2159 287 -2125
rect 229 -2193 241 -2159
rect 275 -2193 287 -2159
rect 229 -2227 287 -2193
rect 229 -2261 241 -2227
rect 275 -2261 287 -2227
rect 229 -2295 287 -2261
rect 229 -2329 241 -2295
rect 275 -2329 287 -2295
rect 229 -2363 287 -2329
rect 229 -2397 241 -2363
rect 275 -2397 287 -2363
rect 229 -2431 287 -2397
rect 229 -2465 241 -2431
rect 275 -2465 287 -2431
rect 229 -2500 287 -2465
rect 487 2465 545 2500
rect 487 2431 499 2465
rect 533 2431 545 2465
rect 487 2397 545 2431
rect 487 2363 499 2397
rect 533 2363 545 2397
rect 487 2329 545 2363
rect 487 2295 499 2329
rect 533 2295 545 2329
rect 487 2261 545 2295
rect 487 2227 499 2261
rect 533 2227 545 2261
rect 487 2193 545 2227
rect 487 2159 499 2193
rect 533 2159 545 2193
rect 487 2125 545 2159
rect 487 2091 499 2125
rect 533 2091 545 2125
rect 487 2057 545 2091
rect 487 2023 499 2057
rect 533 2023 545 2057
rect 487 1989 545 2023
rect 487 1955 499 1989
rect 533 1955 545 1989
rect 487 1921 545 1955
rect 487 1887 499 1921
rect 533 1887 545 1921
rect 487 1853 545 1887
rect 487 1819 499 1853
rect 533 1819 545 1853
rect 487 1785 545 1819
rect 487 1751 499 1785
rect 533 1751 545 1785
rect 487 1717 545 1751
rect 487 1683 499 1717
rect 533 1683 545 1717
rect 487 1649 545 1683
rect 487 1615 499 1649
rect 533 1615 545 1649
rect 487 1581 545 1615
rect 487 1547 499 1581
rect 533 1547 545 1581
rect 487 1513 545 1547
rect 487 1479 499 1513
rect 533 1479 545 1513
rect 487 1445 545 1479
rect 487 1411 499 1445
rect 533 1411 545 1445
rect 487 1377 545 1411
rect 487 1343 499 1377
rect 533 1343 545 1377
rect 487 1309 545 1343
rect 487 1275 499 1309
rect 533 1275 545 1309
rect 487 1241 545 1275
rect 487 1207 499 1241
rect 533 1207 545 1241
rect 487 1173 545 1207
rect 487 1139 499 1173
rect 533 1139 545 1173
rect 487 1105 545 1139
rect 487 1071 499 1105
rect 533 1071 545 1105
rect 487 1037 545 1071
rect 487 1003 499 1037
rect 533 1003 545 1037
rect 487 969 545 1003
rect 487 935 499 969
rect 533 935 545 969
rect 487 901 545 935
rect 487 867 499 901
rect 533 867 545 901
rect 487 833 545 867
rect 487 799 499 833
rect 533 799 545 833
rect 487 765 545 799
rect 487 731 499 765
rect 533 731 545 765
rect 487 697 545 731
rect 487 663 499 697
rect 533 663 545 697
rect 487 629 545 663
rect 487 595 499 629
rect 533 595 545 629
rect 487 561 545 595
rect 487 527 499 561
rect 533 527 545 561
rect 487 493 545 527
rect 487 459 499 493
rect 533 459 545 493
rect 487 425 545 459
rect 487 391 499 425
rect 533 391 545 425
rect 487 357 545 391
rect 487 323 499 357
rect 533 323 545 357
rect 487 289 545 323
rect 487 255 499 289
rect 533 255 545 289
rect 487 221 545 255
rect 487 187 499 221
rect 533 187 545 221
rect 487 153 545 187
rect 487 119 499 153
rect 533 119 545 153
rect 487 85 545 119
rect 487 51 499 85
rect 533 51 545 85
rect 487 17 545 51
rect 487 -17 499 17
rect 533 -17 545 17
rect 487 -51 545 -17
rect 487 -85 499 -51
rect 533 -85 545 -51
rect 487 -119 545 -85
rect 487 -153 499 -119
rect 533 -153 545 -119
rect 487 -187 545 -153
rect 487 -221 499 -187
rect 533 -221 545 -187
rect 487 -255 545 -221
rect 487 -289 499 -255
rect 533 -289 545 -255
rect 487 -323 545 -289
rect 487 -357 499 -323
rect 533 -357 545 -323
rect 487 -391 545 -357
rect 487 -425 499 -391
rect 533 -425 545 -391
rect 487 -459 545 -425
rect 487 -493 499 -459
rect 533 -493 545 -459
rect 487 -527 545 -493
rect 487 -561 499 -527
rect 533 -561 545 -527
rect 487 -595 545 -561
rect 487 -629 499 -595
rect 533 -629 545 -595
rect 487 -663 545 -629
rect 487 -697 499 -663
rect 533 -697 545 -663
rect 487 -731 545 -697
rect 487 -765 499 -731
rect 533 -765 545 -731
rect 487 -799 545 -765
rect 487 -833 499 -799
rect 533 -833 545 -799
rect 487 -867 545 -833
rect 487 -901 499 -867
rect 533 -901 545 -867
rect 487 -935 545 -901
rect 487 -969 499 -935
rect 533 -969 545 -935
rect 487 -1003 545 -969
rect 487 -1037 499 -1003
rect 533 -1037 545 -1003
rect 487 -1071 545 -1037
rect 487 -1105 499 -1071
rect 533 -1105 545 -1071
rect 487 -1139 545 -1105
rect 487 -1173 499 -1139
rect 533 -1173 545 -1139
rect 487 -1207 545 -1173
rect 487 -1241 499 -1207
rect 533 -1241 545 -1207
rect 487 -1275 545 -1241
rect 487 -1309 499 -1275
rect 533 -1309 545 -1275
rect 487 -1343 545 -1309
rect 487 -1377 499 -1343
rect 533 -1377 545 -1343
rect 487 -1411 545 -1377
rect 487 -1445 499 -1411
rect 533 -1445 545 -1411
rect 487 -1479 545 -1445
rect 487 -1513 499 -1479
rect 533 -1513 545 -1479
rect 487 -1547 545 -1513
rect 487 -1581 499 -1547
rect 533 -1581 545 -1547
rect 487 -1615 545 -1581
rect 487 -1649 499 -1615
rect 533 -1649 545 -1615
rect 487 -1683 545 -1649
rect 487 -1717 499 -1683
rect 533 -1717 545 -1683
rect 487 -1751 545 -1717
rect 487 -1785 499 -1751
rect 533 -1785 545 -1751
rect 487 -1819 545 -1785
rect 487 -1853 499 -1819
rect 533 -1853 545 -1819
rect 487 -1887 545 -1853
rect 487 -1921 499 -1887
rect 533 -1921 545 -1887
rect 487 -1955 545 -1921
rect 487 -1989 499 -1955
rect 533 -1989 545 -1955
rect 487 -2023 545 -1989
rect 487 -2057 499 -2023
rect 533 -2057 545 -2023
rect 487 -2091 545 -2057
rect 487 -2125 499 -2091
rect 533 -2125 545 -2091
rect 487 -2159 545 -2125
rect 487 -2193 499 -2159
rect 533 -2193 545 -2159
rect 487 -2227 545 -2193
rect 487 -2261 499 -2227
rect 533 -2261 545 -2227
rect 487 -2295 545 -2261
rect 487 -2329 499 -2295
rect 533 -2329 545 -2295
rect 487 -2363 545 -2329
rect 487 -2397 499 -2363
rect 533 -2397 545 -2363
rect 487 -2431 545 -2397
rect 487 -2465 499 -2431
rect 533 -2465 545 -2431
rect 487 -2500 545 -2465
rect 745 2465 803 2500
rect 745 2431 757 2465
rect 791 2431 803 2465
rect 745 2397 803 2431
rect 745 2363 757 2397
rect 791 2363 803 2397
rect 745 2329 803 2363
rect 745 2295 757 2329
rect 791 2295 803 2329
rect 745 2261 803 2295
rect 745 2227 757 2261
rect 791 2227 803 2261
rect 745 2193 803 2227
rect 745 2159 757 2193
rect 791 2159 803 2193
rect 745 2125 803 2159
rect 745 2091 757 2125
rect 791 2091 803 2125
rect 745 2057 803 2091
rect 745 2023 757 2057
rect 791 2023 803 2057
rect 745 1989 803 2023
rect 745 1955 757 1989
rect 791 1955 803 1989
rect 745 1921 803 1955
rect 745 1887 757 1921
rect 791 1887 803 1921
rect 745 1853 803 1887
rect 745 1819 757 1853
rect 791 1819 803 1853
rect 745 1785 803 1819
rect 745 1751 757 1785
rect 791 1751 803 1785
rect 745 1717 803 1751
rect 745 1683 757 1717
rect 791 1683 803 1717
rect 745 1649 803 1683
rect 745 1615 757 1649
rect 791 1615 803 1649
rect 745 1581 803 1615
rect 745 1547 757 1581
rect 791 1547 803 1581
rect 745 1513 803 1547
rect 745 1479 757 1513
rect 791 1479 803 1513
rect 745 1445 803 1479
rect 745 1411 757 1445
rect 791 1411 803 1445
rect 745 1377 803 1411
rect 745 1343 757 1377
rect 791 1343 803 1377
rect 745 1309 803 1343
rect 745 1275 757 1309
rect 791 1275 803 1309
rect 745 1241 803 1275
rect 745 1207 757 1241
rect 791 1207 803 1241
rect 745 1173 803 1207
rect 745 1139 757 1173
rect 791 1139 803 1173
rect 745 1105 803 1139
rect 745 1071 757 1105
rect 791 1071 803 1105
rect 745 1037 803 1071
rect 745 1003 757 1037
rect 791 1003 803 1037
rect 745 969 803 1003
rect 745 935 757 969
rect 791 935 803 969
rect 745 901 803 935
rect 745 867 757 901
rect 791 867 803 901
rect 745 833 803 867
rect 745 799 757 833
rect 791 799 803 833
rect 745 765 803 799
rect 745 731 757 765
rect 791 731 803 765
rect 745 697 803 731
rect 745 663 757 697
rect 791 663 803 697
rect 745 629 803 663
rect 745 595 757 629
rect 791 595 803 629
rect 745 561 803 595
rect 745 527 757 561
rect 791 527 803 561
rect 745 493 803 527
rect 745 459 757 493
rect 791 459 803 493
rect 745 425 803 459
rect 745 391 757 425
rect 791 391 803 425
rect 745 357 803 391
rect 745 323 757 357
rect 791 323 803 357
rect 745 289 803 323
rect 745 255 757 289
rect 791 255 803 289
rect 745 221 803 255
rect 745 187 757 221
rect 791 187 803 221
rect 745 153 803 187
rect 745 119 757 153
rect 791 119 803 153
rect 745 85 803 119
rect 745 51 757 85
rect 791 51 803 85
rect 745 17 803 51
rect 745 -17 757 17
rect 791 -17 803 17
rect 745 -51 803 -17
rect 745 -85 757 -51
rect 791 -85 803 -51
rect 745 -119 803 -85
rect 745 -153 757 -119
rect 791 -153 803 -119
rect 745 -187 803 -153
rect 745 -221 757 -187
rect 791 -221 803 -187
rect 745 -255 803 -221
rect 745 -289 757 -255
rect 791 -289 803 -255
rect 745 -323 803 -289
rect 745 -357 757 -323
rect 791 -357 803 -323
rect 745 -391 803 -357
rect 745 -425 757 -391
rect 791 -425 803 -391
rect 745 -459 803 -425
rect 745 -493 757 -459
rect 791 -493 803 -459
rect 745 -527 803 -493
rect 745 -561 757 -527
rect 791 -561 803 -527
rect 745 -595 803 -561
rect 745 -629 757 -595
rect 791 -629 803 -595
rect 745 -663 803 -629
rect 745 -697 757 -663
rect 791 -697 803 -663
rect 745 -731 803 -697
rect 745 -765 757 -731
rect 791 -765 803 -731
rect 745 -799 803 -765
rect 745 -833 757 -799
rect 791 -833 803 -799
rect 745 -867 803 -833
rect 745 -901 757 -867
rect 791 -901 803 -867
rect 745 -935 803 -901
rect 745 -969 757 -935
rect 791 -969 803 -935
rect 745 -1003 803 -969
rect 745 -1037 757 -1003
rect 791 -1037 803 -1003
rect 745 -1071 803 -1037
rect 745 -1105 757 -1071
rect 791 -1105 803 -1071
rect 745 -1139 803 -1105
rect 745 -1173 757 -1139
rect 791 -1173 803 -1139
rect 745 -1207 803 -1173
rect 745 -1241 757 -1207
rect 791 -1241 803 -1207
rect 745 -1275 803 -1241
rect 745 -1309 757 -1275
rect 791 -1309 803 -1275
rect 745 -1343 803 -1309
rect 745 -1377 757 -1343
rect 791 -1377 803 -1343
rect 745 -1411 803 -1377
rect 745 -1445 757 -1411
rect 791 -1445 803 -1411
rect 745 -1479 803 -1445
rect 745 -1513 757 -1479
rect 791 -1513 803 -1479
rect 745 -1547 803 -1513
rect 745 -1581 757 -1547
rect 791 -1581 803 -1547
rect 745 -1615 803 -1581
rect 745 -1649 757 -1615
rect 791 -1649 803 -1615
rect 745 -1683 803 -1649
rect 745 -1717 757 -1683
rect 791 -1717 803 -1683
rect 745 -1751 803 -1717
rect 745 -1785 757 -1751
rect 791 -1785 803 -1751
rect 745 -1819 803 -1785
rect 745 -1853 757 -1819
rect 791 -1853 803 -1819
rect 745 -1887 803 -1853
rect 745 -1921 757 -1887
rect 791 -1921 803 -1887
rect 745 -1955 803 -1921
rect 745 -1989 757 -1955
rect 791 -1989 803 -1955
rect 745 -2023 803 -1989
rect 745 -2057 757 -2023
rect 791 -2057 803 -2023
rect 745 -2091 803 -2057
rect 745 -2125 757 -2091
rect 791 -2125 803 -2091
rect 745 -2159 803 -2125
rect 745 -2193 757 -2159
rect 791 -2193 803 -2159
rect 745 -2227 803 -2193
rect 745 -2261 757 -2227
rect 791 -2261 803 -2227
rect 745 -2295 803 -2261
rect 745 -2329 757 -2295
rect 791 -2329 803 -2295
rect 745 -2363 803 -2329
rect 745 -2397 757 -2363
rect 791 -2397 803 -2363
rect 745 -2431 803 -2397
rect 745 -2465 757 -2431
rect 791 -2465 803 -2431
rect 745 -2500 803 -2465
rect 1003 2465 1061 2500
rect 1003 2431 1015 2465
rect 1049 2431 1061 2465
rect 1003 2397 1061 2431
rect 1003 2363 1015 2397
rect 1049 2363 1061 2397
rect 1003 2329 1061 2363
rect 1003 2295 1015 2329
rect 1049 2295 1061 2329
rect 1003 2261 1061 2295
rect 1003 2227 1015 2261
rect 1049 2227 1061 2261
rect 1003 2193 1061 2227
rect 1003 2159 1015 2193
rect 1049 2159 1061 2193
rect 1003 2125 1061 2159
rect 1003 2091 1015 2125
rect 1049 2091 1061 2125
rect 1003 2057 1061 2091
rect 1003 2023 1015 2057
rect 1049 2023 1061 2057
rect 1003 1989 1061 2023
rect 1003 1955 1015 1989
rect 1049 1955 1061 1989
rect 1003 1921 1061 1955
rect 1003 1887 1015 1921
rect 1049 1887 1061 1921
rect 1003 1853 1061 1887
rect 1003 1819 1015 1853
rect 1049 1819 1061 1853
rect 1003 1785 1061 1819
rect 1003 1751 1015 1785
rect 1049 1751 1061 1785
rect 1003 1717 1061 1751
rect 1003 1683 1015 1717
rect 1049 1683 1061 1717
rect 1003 1649 1061 1683
rect 1003 1615 1015 1649
rect 1049 1615 1061 1649
rect 1003 1581 1061 1615
rect 1003 1547 1015 1581
rect 1049 1547 1061 1581
rect 1003 1513 1061 1547
rect 1003 1479 1015 1513
rect 1049 1479 1061 1513
rect 1003 1445 1061 1479
rect 1003 1411 1015 1445
rect 1049 1411 1061 1445
rect 1003 1377 1061 1411
rect 1003 1343 1015 1377
rect 1049 1343 1061 1377
rect 1003 1309 1061 1343
rect 1003 1275 1015 1309
rect 1049 1275 1061 1309
rect 1003 1241 1061 1275
rect 1003 1207 1015 1241
rect 1049 1207 1061 1241
rect 1003 1173 1061 1207
rect 1003 1139 1015 1173
rect 1049 1139 1061 1173
rect 1003 1105 1061 1139
rect 1003 1071 1015 1105
rect 1049 1071 1061 1105
rect 1003 1037 1061 1071
rect 1003 1003 1015 1037
rect 1049 1003 1061 1037
rect 1003 969 1061 1003
rect 1003 935 1015 969
rect 1049 935 1061 969
rect 1003 901 1061 935
rect 1003 867 1015 901
rect 1049 867 1061 901
rect 1003 833 1061 867
rect 1003 799 1015 833
rect 1049 799 1061 833
rect 1003 765 1061 799
rect 1003 731 1015 765
rect 1049 731 1061 765
rect 1003 697 1061 731
rect 1003 663 1015 697
rect 1049 663 1061 697
rect 1003 629 1061 663
rect 1003 595 1015 629
rect 1049 595 1061 629
rect 1003 561 1061 595
rect 1003 527 1015 561
rect 1049 527 1061 561
rect 1003 493 1061 527
rect 1003 459 1015 493
rect 1049 459 1061 493
rect 1003 425 1061 459
rect 1003 391 1015 425
rect 1049 391 1061 425
rect 1003 357 1061 391
rect 1003 323 1015 357
rect 1049 323 1061 357
rect 1003 289 1061 323
rect 1003 255 1015 289
rect 1049 255 1061 289
rect 1003 221 1061 255
rect 1003 187 1015 221
rect 1049 187 1061 221
rect 1003 153 1061 187
rect 1003 119 1015 153
rect 1049 119 1061 153
rect 1003 85 1061 119
rect 1003 51 1015 85
rect 1049 51 1061 85
rect 1003 17 1061 51
rect 1003 -17 1015 17
rect 1049 -17 1061 17
rect 1003 -51 1061 -17
rect 1003 -85 1015 -51
rect 1049 -85 1061 -51
rect 1003 -119 1061 -85
rect 1003 -153 1015 -119
rect 1049 -153 1061 -119
rect 1003 -187 1061 -153
rect 1003 -221 1015 -187
rect 1049 -221 1061 -187
rect 1003 -255 1061 -221
rect 1003 -289 1015 -255
rect 1049 -289 1061 -255
rect 1003 -323 1061 -289
rect 1003 -357 1015 -323
rect 1049 -357 1061 -323
rect 1003 -391 1061 -357
rect 1003 -425 1015 -391
rect 1049 -425 1061 -391
rect 1003 -459 1061 -425
rect 1003 -493 1015 -459
rect 1049 -493 1061 -459
rect 1003 -527 1061 -493
rect 1003 -561 1015 -527
rect 1049 -561 1061 -527
rect 1003 -595 1061 -561
rect 1003 -629 1015 -595
rect 1049 -629 1061 -595
rect 1003 -663 1061 -629
rect 1003 -697 1015 -663
rect 1049 -697 1061 -663
rect 1003 -731 1061 -697
rect 1003 -765 1015 -731
rect 1049 -765 1061 -731
rect 1003 -799 1061 -765
rect 1003 -833 1015 -799
rect 1049 -833 1061 -799
rect 1003 -867 1061 -833
rect 1003 -901 1015 -867
rect 1049 -901 1061 -867
rect 1003 -935 1061 -901
rect 1003 -969 1015 -935
rect 1049 -969 1061 -935
rect 1003 -1003 1061 -969
rect 1003 -1037 1015 -1003
rect 1049 -1037 1061 -1003
rect 1003 -1071 1061 -1037
rect 1003 -1105 1015 -1071
rect 1049 -1105 1061 -1071
rect 1003 -1139 1061 -1105
rect 1003 -1173 1015 -1139
rect 1049 -1173 1061 -1139
rect 1003 -1207 1061 -1173
rect 1003 -1241 1015 -1207
rect 1049 -1241 1061 -1207
rect 1003 -1275 1061 -1241
rect 1003 -1309 1015 -1275
rect 1049 -1309 1061 -1275
rect 1003 -1343 1061 -1309
rect 1003 -1377 1015 -1343
rect 1049 -1377 1061 -1343
rect 1003 -1411 1061 -1377
rect 1003 -1445 1015 -1411
rect 1049 -1445 1061 -1411
rect 1003 -1479 1061 -1445
rect 1003 -1513 1015 -1479
rect 1049 -1513 1061 -1479
rect 1003 -1547 1061 -1513
rect 1003 -1581 1015 -1547
rect 1049 -1581 1061 -1547
rect 1003 -1615 1061 -1581
rect 1003 -1649 1015 -1615
rect 1049 -1649 1061 -1615
rect 1003 -1683 1061 -1649
rect 1003 -1717 1015 -1683
rect 1049 -1717 1061 -1683
rect 1003 -1751 1061 -1717
rect 1003 -1785 1015 -1751
rect 1049 -1785 1061 -1751
rect 1003 -1819 1061 -1785
rect 1003 -1853 1015 -1819
rect 1049 -1853 1061 -1819
rect 1003 -1887 1061 -1853
rect 1003 -1921 1015 -1887
rect 1049 -1921 1061 -1887
rect 1003 -1955 1061 -1921
rect 1003 -1989 1015 -1955
rect 1049 -1989 1061 -1955
rect 1003 -2023 1061 -1989
rect 1003 -2057 1015 -2023
rect 1049 -2057 1061 -2023
rect 1003 -2091 1061 -2057
rect 1003 -2125 1015 -2091
rect 1049 -2125 1061 -2091
rect 1003 -2159 1061 -2125
rect 1003 -2193 1015 -2159
rect 1049 -2193 1061 -2159
rect 1003 -2227 1061 -2193
rect 1003 -2261 1015 -2227
rect 1049 -2261 1061 -2227
rect 1003 -2295 1061 -2261
rect 1003 -2329 1015 -2295
rect 1049 -2329 1061 -2295
rect 1003 -2363 1061 -2329
rect 1003 -2397 1015 -2363
rect 1049 -2397 1061 -2363
rect 1003 -2431 1061 -2397
rect 1003 -2465 1015 -2431
rect 1049 -2465 1061 -2431
rect 1003 -2500 1061 -2465
rect 1261 2465 1319 2500
rect 1261 2431 1273 2465
rect 1307 2431 1319 2465
rect 1261 2397 1319 2431
rect 1261 2363 1273 2397
rect 1307 2363 1319 2397
rect 1261 2329 1319 2363
rect 1261 2295 1273 2329
rect 1307 2295 1319 2329
rect 1261 2261 1319 2295
rect 1261 2227 1273 2261
rect 1307 2227 1319 2261
rect 1261 2193 1319 2227
rect 1261 2159 1273 2193
rect 1307 2159 1319 2193
rect 1261 2125 1319 2159
rect 1261 2091 1273 2125
rect 1307 2091 1319 2125
rect 1261 2057 1319 2091
rect 1261 2023 1273 2057
rect 1307 2023 1319 2057
rect 1261 1989 1319 2023
rect 1261 1955 1273 1989
rect 1307 1955 1319 1989
rect 1261 1921 1319 1955
rect 1261 1887 1273 1921
rect 1307 1887 1319 1921
rect 1261 1853 1319 1887
rect 1261 1819 1273 1853
rect 1307 1819 1319 1853
rect 1261 1785 1319 1819
rect 1261 1751 1273 1785
rect 1307 1751 1319 1785
rect 1261 1717 1319 1751
rect 1261 1683 1273 1717
rect 1307 1683 1319 1717
rect 1261 1649 1319 1683
rect 1261 1615 1273 1649
rect 1307 1615 1319 1649
rect 1261 1581 1319 1615
rect 1261 1547 1273 1581
rect 1307 1547 1319 1581
rect 1261 1513 1319 1547
rect 1261 1479 1273 1513
rect 1307 1479 1319 1513
rect 1261 1445 1319 1479
rect 1261 1411 1273 1445
rect 1307 1411 1319 1445
rect 1261 1377 1319 1411
rect 1261 1343 1273 1377
rect 1307 1343 1319 1377
rect 1261 1309 1319 1343
rect 1261 1275 1273 1309
rect 1307 1275 1319 1309
rect 1261 1241 1319 1275
rect 1261 1207 1273 1241
rect 1307 1207 1319 1241
rect 1261 1173 1319 1207
rect 1261 1139 1273 1173
rect 1307 1139 1319 1173
rect 1261 1105 1319 1139
rect 1261 1071 1273 1105
rect 1307 1071 1319 1105
rect 1261 1037 1319 1071
rect 1261 1003 1273 1037
rect 1307 1003 1319 1037
rect 1261 969 1319 1003
rect 1261 935 1273 969
rect 1307 935 1319 969
rect 1261 901 1319 935
rect 1261 867 1273 901
rect 1307 867 1319 901
rect 1261 833 1319 867
rect 1261 799 1273 833
rect 1307 799 1319 833
rect 1261 765 1319 799
rect 1261 731 1273 765
rect 1307 731 1319 765
rect 1261 697 1319 731
rect 1261 663 1273 697
rect 1307 663 1319 697
rect 1261 629 1319 663
rect 1261 595 1273 629
rect 1307 595 1319 629
rect 1261 561 1319 595
rect 1261 527 1273 561
rect 1307 527 1319 561
rect 1261 493 1319 527
rect 1261 459 1273 493
rect 1307 459 1319 493
rect 1261 425 1319 459
rect 1261 391 1273 425
rect 1307 391 1319 425
rect 1261 357 1319 391
rect 1261 323 1273 357
rect 1307 323 1319 357
rect 1261 289 1319 323
rect 1261 255 1273 289
rect 1307 255 1319 289
rect 1261 221 1319 255
rect 1261 187 1273 221
rect 1307 187 1319 221
rect 1261 153 1319 187
rect 1261 119 1273 153
rect 1307 119 1319 153
rect 1261 85 1319 119
rect 1261 51 1273 85
rect 1307 51 1319 85
rect 1261 17 1319 51
rect 1261 -17 1273 17
rect 1307 -17 1319 17
rect 1261 -51 1319 -17
rect 1261 -85 1273 -51
rect 1307 -85 1319 -51
rect 1261 -119 1319 -85
rect 1261 -153 1273 -119
rect 1307 -153 1319 -119
rect 1261 -187 1319 -153
rect 1261 -221 1273 -187
rect 1307 -221 1319 -187
rect 1261 -255 1319 -221
rect 1261 -289 1273 -255
rect 1307 -289 1319 -255
rect 1261 -323 1319 -289
rect 1261 -357 1273 -323
rect 1307 -357 1319 -323
rect 1261 -391 1319 -357
rect 1261 -425 1273 -391
rect 1307 -425 1319 -391
rect 1261 -459 1319 -425
rect 1261 -493 1273 -459
rect 1307 -493 1319 -459
rect 1261 -527 1319 -493
rect 1261 -561 1273 -527
rect 1307 -561 1319 -527
rect 1261 -595 1319 -561
rect 1261 -629 1273 -595
rect 1307 -629 1319 -595
rect 1261 -663 1319 -629
rect 1261 -697 1273 -663
rect 1307 -697 1319 -663
rect 1261 -731 1319 -697
rect 1261 -765 1273 -731
rect 1307 -765 1319 -731
rect 1261 -799 1319 -765
rect 1261 -833 1273 -799
rect 1307 -833 1319 -799
rect 1261 -867 1319 -833
rect 1261 -901 1273 -867
rect 1307 -901 1319 -867
rect 1261 -935 1319 -901
rect 1261 -969 1273 -935
rect 1307 -969 1319 -935
rect 1261 -1003 1319 -969
rect 1261 -1037 1273 -1003
rect 1307 -1037 1319 -1003
rect 1261 -1071 1319 -1037
rect 1261 -1105 1273 -1071
rect 1307 -1105 1319 -1071
rect 1261 -1139 1319 -1105
rect 1261 -1173 1273 -1139
rect 1307 -1173 1319 -1139
rect 1261 -1207 1319 -1173
rect 1261 -1241 1273 -1207
rect 1307 -1241 1319 -1207
rect 1261 -1275 1319 -1241
rect 1261 -1309 1273 -1275
rect 1307 -1309 1319 -1275
rect 1261 -1343 1319 -1309
rect 1261 -1377 1273 -1343
rect 1307 -1377 1319 -1343
rect 1261 -1411 1319 -1377
rect 1261 -1445 1273 -1411
rect 1307 -1445 1319 -1411
rect 1261 -1479 1319 -1445
rect 1261 -1513 1273 -1479
rect 1307 -1513 1319 -1479
rect 1261 -1547 1319 -1513
rect 1261 -1581 1273 -1547
rect 1307 -1581 1319 -1547
rect 1261 -1615 1319 -1581
rect 1261 -1649 1273 -1615
rect 1307 -1649 1319 -1615
rect 1261 -1683 1319 -1649
rect 1261 -1717 1273 -1683
rect 1307 -1717 1319 -1683
rect 1261 -1751 1319 -1717
rect 1261 -1785 1273 -1751
rect 1307 -1785 1319 -1751
rect 1261 -1819 1319 -1785
rect 1261 -1853 1273 -1819
rect 1307 -1853 1319 -1819
rect 1261 -1887 1319 -1853
rect 1261 -1921 1273 -1887
rect 1307 -1921 1319 -1887
rect 1261 -1955 1319 -1921
rect 1261 -1989 1273 -1955
rect 1307 -1989 1319 -1955
rect 1261 -2023 1319 -1989
rect 1261 -2057 1273 -2023
rect 1307 -2057 1319 -2023
rect 1261 -2091 1319 -2057
rect 1261 -2125 1273 -2091
rect 1307 -2125 1319 -2091
rect 1261 -2159 1319 -2125
rect 1261 -2193 1273 -2159
rect 1307 -2193 1319 -2159
rect 1261 -2227 1319 -2193
rect 1261 -2261 1273 -2227
rect 1307 -2261 1319 -2227
rect 1261 -2295 1319 -2261
rect 1261 -2329 1273 -2295
rect 1307 -2329 1319 -2295
rect 1261 -2363 1319 -2329
rect 1261 -2397 1273 -2363
rect 1307 -2397 1319 -2363
rect 1261 -2431 1319 -2397
rect 1261 -2465 1273 -2431
rect 1307 -2465 1319 -2431
rect 1261 -2500 1319 -2465
<< ndiffc >>
rect -1307 2431 -1273 2465
rect -1307 2363 -1273 2397
rect -1307 2295 -1273 2329
rect -1307 2227 -1273 2261
rect -1307 2159 -1273 2193
rect -1307 2091 -1273 2125
rect -1307 2023 -1273 2057
rect -1307 1955 -1273 1989
rect -1307 1887 -1273 1921
rect -1307 1819 -1273 1853
rect -1307 1751 -1273 1785
rect -1307 1683 -1273 1717
rect -1307 1615 -1273 1649
rect -1307 1547 -1273 1581
rect -1307 1479 -1273 1513
rect -1307 1411 -1273 1445
rect -1307 1343 -1273 1377
rect -1307 1275 -1273 1309
rect -1307 1207 -1273 1241
rect -1307 1139 -1273 1173
rect -1307 1071 -1273 1105
rect -1307 1003 -1273 1037
rect -1307 935 -1273 969
rect -1307 867 -1273 901
rect -1307 799 -1273 833
rect -1307 731 -1273 765
rect -1307 663 -1273 697
rect -1307 595 -1273 629
rect -1307 527 -1273 561
rect -1307 459 -1273 493
rect -1307 391 -1273 425
rect -1307 323 -1273 357
rect -1307 255 -1273 289
rect -1307 187 -1273 221
rect -1307 119 -1273 153
rect -1307 51 -1273 85
rect -1307 -17 -1273 17
rect -1307 -85 -1273 -51
rect -1307 -153 -1273 -119
rect -1307 -221 -1273 -187
rect -1307 -289 -1273 -255
rect -1307 -357 -1273 -323
rect -1307 -425 -1273 -391
rect -1307 -493 -1273 -459
rect -1307 -561 -1273 -527
rect -1307 -629 -1273 -595
rect -1307 -697 -1273 -663
rect -1307 -765 -1273 -731
rect -1307 -833 -1273 -799
rect -1307 -901 -1273 -867
rect -1307 -969 -1273 -935
rect -1307 -1037 -1273 -1003
rect -1307 -1105 -1273 -1071
rect -1307 -1173 -1273 -1139
rect -1307 -1241 -1273 -1207
rect -1307 -1309 -1273 -1275
rect -1307 -1377 -1273 -1343
rect -1307 -1445 -1273 -1411
rect -1307 -1513 -1273 -1479
rect -1307 -1581 -1273 -1547
rect -1307 -1649 -1273 -1615
rect -1307 -1717 -1273 -1683
rect -1307 -1785 -1273 -1751
rect -1307 -1853 -1273 -1819
rect -1307 -1921 -1273 -1887
rect -1307 -1989 -1273 -1955
rect -1307 -2057 -1273 -2023
rect -1307 -2125 -1273 -2091
rect -1307 -2193 -1273 -2159
rect -1307 -2261 -1273 -2227
rect -1307 -2329 -1273 -2295
rect -1307 -2397 -1273 -2363
rect -1307 -2465 -1273 -2431
rect -1049 2431 -1015 2465
rect -1049 2363 -1015 2397
rect -1049 2295 -1015 2329
rect -1049 2227 -1015 2261
rect -1049 2159 -1015 2193
rect -1049 2091 -1015 2125
rect -1049 2023 -1015 2057
rect -1049 1955 -1015 1989
rect -1049 1887 -1015 1921
rect -1049 1819 -1015 1853
rect -1049 1751 -1015 1785
rect -1049 1683 -1015 1717
rect -1049 1615 -1015 1649
rect -1049 1547 -1015 1581
rect -1049 1479 -1015 1513
rect -1049 1411 -1015 1445
rect -1049 1343 -1015 1377
rect -1049 1275 -1015 1309
rect -1049 1207 -1015 1241
rect -1049 1139 -1015 1173
rect -1049 1071 -1015 1105
rect -1049 1003 -1015 1037
rect -1049 935 -1015 969
rect -1049 867 -1015 901
rect -1049 799 -1015 833
rect -1049 731 -1015 765
rect -1049 663 -1015 697
rect -1049 595 -1015 629
rect -1049 527 -1015 561
rect -1049 459 -1015 493
rect -1049 391 -1015 425
rect -1049 323 -1015 357
rect -1049 255 -1015 289
rect -1049 187 -1015 221
rect -1049 119 -1015 153
rect -1049 51 -1015 85
rect -1049 -17 -1015 17
rect -1049 -85 -1015 -51
rect -1049 -153 -1015 -119
rect -1049 -221 -1015 -187
rect -1049 -289 -1015 -255
rect -1049 -357 -1015 -323
rect -1049 -425 -1015 -391
rect -1049 -493 -1015 -459
rect -1049 -561 -1015 -527
rect -1049 -629 -1015 -595
rect -1049 -697 -1015 -663
rect -1049 -765 -1015 -731
rect -1049 -833 -1015 -799
rect -1049 -901 -1015 -867
rect -1049 -969 -1015 -935
rect -1049 -1037 -1015 -1003
rect -1049 -1105 -1015 -1071
rect -1049 -1173 -1015 -1139
rect -1049 -1241 -1015 -1207
rect -1049 -1309 -1015 -1275
rect -1049 -1377 -1015 -1343
rect -1049 -1445 -1015 -1411
rect -1049 -1513 -1015 -1479
rect -1049 -1581 -1015 -1547
rect -1049 -1649 -1015 -1615
rect -1049 -1717 -1015 -1683
rect -1049 -1785 -1015 -1751
rect -1049 -1853 -1015 -1819
rect -1049 -1921 -1015 -1887
rect -1049 -1989 -1015 -1955
rect -1049 -2057 -1015 -2023
rect -1049 -2125 -1015 -2091
rect -1049 -2193 -1015 -2159
rect -1049 -2261 -1015 -2227
rect -1049 -2329 -1015 -2295
rect -1049 -2397 -1015 -2363
rect -1049 -2465 -1015 -2431
rect -791 2431 -757 2465
rect -791 2363 -757 2397
rect -791 2295 -757 2329
rect -791 2227 -757 2261
rect -791 2159 -757 2193
rect -791 2091 -757 2125
rect -791 2023 -757 2057
rect -791 1955 -757 1989
rect -791 1887 -757 1921
rect -791 1819 -757 1853
rect -791 1751 -757 1785
rect -791 1683 -757 1717
rect -791 1615 -757 1649
rect -791 1547 -757 1581
rect -791 1479 -757 1513
rect -791 1411 -757 1445
rect -791 1343 -757 1377
rect -791 1275 -757 1309
rect -791 1207 -757 1241
rect -791 1139 -757 1173
rect -791 1071 -757 1105
rect -791 1003 -757 1037
rect -791 935 -757 969
rect -791 867 -757 901
rect -791 799 -757 833
rect -791 731 -757 765
rect -791 663 -757 697
rect -791 595 -757 629
rect -791 527 -757 561
rect -791 459 -757 493
rect -791 391 -757 425
rect -791 323 -757 357
rect -791 255 -757 289
rect -791 187 -757 221
rect -791 119 -757 153
rect -791 51 -757 85
rect -791 -17 -757 17
rect -791 -85 -757 -51
rect -791 -153 -757 -119
rect -791 -221 -757 -187
rect -791 -289 -757 -255
rect -791 -357 -757 -323
rect -791 -425 -757 -391
rect -791 -493 -757 -459
rect -791 -561 -757 -527
rect -791 -629 -757 -595
rect -791 -697 -757 -663
rect -791 -765 -757 -731
rect -791 -833 -757 -799
rect -791 -901 -757 -867
rect -791 -969 -757 -935
rect -791 -1037 -757 -1003
rect -791 -1105 -757 -1071
rect -791 -1173 -757 -1139
rect -791 -1241 -757 -1207
rect -791 -1309 -757 -1275
rect -791 -1377 -757 -1343
rect -791 -1445 -757 -1411
rect -791 -1513 -757 -1479
rect -791 -1581 -757 -1547
rect -791 -1649 -757 -1615
rect -791 -1717 -757 -1683
rect -791 -1785 -757 -1751
rect -791 -1853 -757 -1819
rect -791 -1921 -757 -1887
rect -791 -1989 -757 -1955
rect -791 -2057 -757 -2023
rect -791 -2125 -757 -2091
rect -791 -2193 -757 -2159
rect -791 -2261 -757 -2227
rect -791 -2329 -757 -2295
rect -791 -2397 -757 -2363
rect -791 -2465 -757 -2431
rect -533 2431 -499 2465
rect -533 2363 -499 2397
rect -533 2295 -499 2329
rect -533 2227 -499 2261
rect -533 2159 -499 2193
rect -533 2091 -499 2125
rect -533 2023 -499 2057
rect -533 1955 -499 1989
rect -533 1887 -499 1921
rect -533 1819 -499 1853
rect -533 1751 -499 1785
rect -533 1683 -499 1717
rect -533 1615 -499 1649
rect -533 1547 -499 1581
rect -533 1479 -499 1513
rect -533 1411 -499 1445
rect -533 1343 -499 1377
rect -533 1275 -499 1309
rect -533 1207 -499 1241
rect -533 1139 -499 1173
rect -533 1071 -499 1105
rect -533 1003 -499 1037
rect -533 935 -499 969
rect -533 867 -499 901
rect -533 799 -499 833
rect -533 731 -499 765
rect -533 663 -499 697
rect -533 595 -499 629
rect -533 527 -499 561
rect -533 459 -499 493
rect -533 391 -499 425
rect -533 323 -499 357
rect -533 255 -499 289
rect -533 187 -499 221
rect -533 119 -499 153
rect -533 51 -499 85
rect -533 -17 -499 17
rect -533 -85 -499 -51
rect -533 -153 -499 -119
rect -533 -221 -499 -187
rect -533 -289 -499 -255
rect -533 -357 -499 -323
rect -533 -425 -499 -391
rect -533 -493 -499 -459
rect -533 -561 -499 -527
rect -533 -629 -499 -595
rect -533 -697 -499 -663
rect -533 -765 -499 -731
rect -533 -833 -499 -799
rect -533 -901 -499 -867
rect -533 -969 -499 -935
rect -533 -1037 -499 -1003
rect -533 -1105 -499 -1071
rect -533 -1173 -499 -1139
rect -533 -1241 -499 -1207
rect -533 -1309 -499 -1275
rect -533 -1377 -499 -1343
rect -533 -1445 -499 -1411
rect -533 -1513 -499 -1479
rect -533 -1581 -499 -1547
rect -533 -1649 -499 -1615
rect -533 -1717 -499 -1683
rect -533 -1785 -499 -1751
rect -533 -1853 -499 -1819
rect -533 -1921 -499 -1887
rect -533 -1989 -499 -1955
rect -533 -2057 -499 -2023
rect -533 -2125 -499 -2091
rect -533 -2193 -499 -2159
rect -533 -2261 -499 -2227
rect -533 -2329 -499 -2295
rect -533 -2397 -499 -2363
rect -533 -2465 -499 -2431
rect -275 2431 -241 2465
rect -275 2363 -241 2397
rect -275 2295 -241 2329
rect -275 2227 -241 2261
rect -275 2159 -241 2193
rect -275 2091 -241 2125
rect -275 2023 -241 2057
rect -275 1955 -241 1989
rect -275 1887 -241 1921
rect -275 1819 -241 1853
rect -275 1751 -241 1785
rect -275 1683 -241 1717
rect -275 1615 -241 1649
rect -275 1547 -241 1581
rect -275 1479 -241 1513
rect -275 1411 -241 1445
rect -275 1343 -241 1377
rect -275 1275 -241 1309
rect -275 1207 -241 1241
rect -275 1139 -241 1173
rect -275 1071 -241 1105
rect -275 1003 -241 1037
rect -275 935 -241 969
rect -275 867 -241 901
rect -275 799 -241 833
rect -275 731 -241 765
rect -275 663 -241 697
rect -275 595 -241 629
rect -275 527 -241 561
rect -275 459 -241 493
rect -275 391 -241 425
rect -275 323 -241 357
rect -275 255 -241 289
rect -275 187 -241 221
rect -275 119 -241 153
rect -275 51 -241 85
rect -275 -17 -241 17
rect -275 -85 -241 -51
rect -275 -153 -241 -119
rect -275 -221 -241 -187
rect -275 -289 -241 -255
rect -275 -357 -241 -323
rect -275 -425 -241 -391
rect -275 -493 -241 -459
rect -275 -561 -241 -527
rect -275 -629 -241 -595
rect -275 -697 -241 -663
rect -275 -765 -241 -731
rect -275 -833 -241 -799
rect -275 -901 -241 -867
rect -275 -969 -241 -935
rect -275 -1037 -241 -1003
rect -275 -1105 -241 -1071
rect -275 -1173 -241 -1139
rect -275 -1241 -241 -1207
rect -275 -1309 -241 -1275
rect -275 -1377 -241 -1343
rect -275 -1445 -241 -1411
rect -275 -1513 -241 -1479
rect -275 -1581 -241 -1547
rect -275 -1649 -241 -1615
rect -275 -1717 -241 -1683
rect -275 -1785 -241 -1751
rect -275 -1853 -241 -1819
rect -275 -1921 -241 -1887
rect -275 -1989 -241 -1955
rect -275 -2057 -241 -2023
rect -275 -2125 -241 -2091
rect -275 -2193 -241 -2159
rect -275 -2261 -241 -2227
rect -275 -2329 -241 -2295
rect -275 -2397 -241 -2363
rect -275 -2465 -241 -2431
rect -17 2431 17 2465
rect -17 2363 17 2397
rect -17 2295 17 2329
rect -17 2227 17 2261
rect -17 2159 17 2193
rect -17 2091 17 2125
rect -17 2023 17 2057
rect -17 1955 17 1989
rect -17 1887 17 1921
rect -17 1819 17 1853
rect -17 1751 17 1785
rect -17 1683 17 1717
rect -17 1615 17 1649
rect -17 1547 17 1581
rect -17 1479 17 1513
rect -17 1411 17 1445
rect -17 1343 17 1377
rect -17 1275 17 1309
rect -17 1207 17 1241
rect -17 1139 17 1173
rect -17 1071 17 1105
rect -17 1003 17 1037
rect -17 935 17 969
rect -17 867 17 901
rect -17 799 17 833
rect -17 731 17 765
rect -17 663 17 697
rect -17 595 17 629
rect -17 527 17 561
rect -17 459 17 493
rect -17 391 17 425
rect -17 323 17 357
rect -17 255 17 289
rect -17 187 17 221
rect -17 119 17 153
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect -17 -153 17 -119
rect -17 -221 17 -187
rect -17 -289 17 -255
rect -17 -357 17 -323
rect -17 -425 17 -391
rect -17 -493 17 -459
rect -17 -561 17 -527
rect -17 -629 17 -595
rect -17 -697 17 -663
rect -17 -765 17 -731
rect -17 -833 17 -799
rect -17 -901 17 -867
rect -17 -969 17 -935
rect -17 -1037 17 -1003
rect -17 -1105 17 -1071
rect -17 -1173 17 -1139
rect -17 -1241 17 -1207
rect -17 -1309 17 -1275
rect -17 -1377 17 -1343
rect -17 -1445 17 -1411
rect -17 -1513 17 -1479
rect -17 -1581 17 -1547
rect -17 -1649 17 -1615
rect -17 -1717 17 -1683
rect -17 -1785 17 -1751
rect -17 -1853 17 -1819
rect -17 -1921 17 -1887
rect -17 -1989 17 -1955
rect -17 -2057 17 -2023
rect -17 -2125 17 -2091
rect -17 -2193 17 -2159
rect -17 -2261 17 -2227
rect -17 -2329 17 -2295
rect -17 -2397 17 -2363
rect -17 -2465 17 -2431
rect 241 2431 275 2465
rect 241 2363 275 2397
rect 241 2295 275 2329
rect 241 2227 275 2261
rect 241 2159 275 2193
rect 241 2091 275 2125
rect 241 2023 275 2057
rect 241 1955 275 1989
rect 241 1887 275 1921
rect 241 1819 275 1853
rect 241 1751 275 1785
rect 241 1683 275 1717
rect 241 1615 275 1649
rect 241 1547 275 1581
rect 241 1479 275 1513
rect 241 1411 275 1445
rect 241 1343 275 1377
rect 241 1275 275 1309
rect 241 1207 275 1241
rect 241 1139 275 1173
rect 241 1071 275 1105
rect 241 1003 275 1037
rect 241 935 275 969
rect 241 867 275 901
rect 241 799 275 833
rect 241 731 275 765
rect 241 663 275 697
rect 241 595 275 629
rect 241 527 275 561
rect 241 459 275 493
rect 241 391 275 425
rect 241 323 275 357
rect 241 255 275 289
rect 241 187 275 221
rect 241 119 275 153
rect 241 51 275 85
rect 241 -17 275 17
rect 241 -85 275 -51
rect 241 -153 275 -119
rect 241 -221 275 -187
rect 241 -289 275 -255
rect 241 -357 275 -323
rect 241 -425 275 -391
rect 241 -493 275 -459
rect 241 -561 275 -527
rect 241 -629 275 -595
rect 241 -697 275 -663
rect 241 -765 275 -731
rect 241 -833 275 -799
rect 241 -901 275 -867
rect 241 -969 275 -935
rect 241 -1037 275 -1003
rect 241 -1105 275 -1071
rect 241 -1173 275 -1139
rect 241 -1241 275 -1207
rect 241 -1309 275 -1275
rect 241 -1377 275 -1343
rect 241 -1445 275 -1411
rect 241 -1513 275 -1479
rect 241 -1581 275 -1547
rect 241 -1649 275 -1615
rect 241 -1717 275 -1683
rect 241 -1785 275 -1751
rect 241 -1853 275 -1819
rect 241 -1921 275 -1887
rect 241 -1989 275 -1955
rect 241 -2057 275 -2023
rect 241 -2125 275 -2091
rect 241 -2193 275 -2159
rect 241 -2261 275 -2227
rect 241 -2329 275 -2295
rect 241 -2397 275 -2363
rect 241 -2465 275 -2431
rect 499 2431 533 2465
rect 499 2363 533 2397
rect 499 2295 533 2329
rect 499 2227 533 2261
rect 499 2159 533 2193
rect 499 2091 533 2125
rect 499 2023 533 2057
rect 499 1955 533 1989
rect 499 1887 533 1921
rect 499 1819 533 1853
rect 499 1751 533 1785
rect 499 1683 533 1717
rect 499 1615 533 1649
rect 499 1547 533 1581
rect 499 1479 533 1513
rect 499 1411 533 1445
rect 499 1343 533 1377
rect 499 1275 533 1309
rect 499 1207 533 1241
rect 499 1139 533 1173
rect 499 1071 533 1105
rect 499 1003 533 1037
rect 499 935 533 969
rect 499 867 533 901
rect 499 799 533 833
rect 499 731 533 765
rect 499 663 533 697
rect 499 595 533 629
rect 499 527 533 561
rect 499 459 533 493
rect 499 391 533 425
rect 499 323 533 357
rect 499 255 533 289
rect 499 187 533 221
rect 499 119 533 153
rect 499 51 533 85
rect 499 -17 533 17
rect 499 -85 533 -51
rect 499 -153 533 -119
rect 499 -221 533 -187
rect 499 -289 533 -255
rect 499 -357 533 -323
rect 499 -425 533 -391
rect 499 -493 533 -459
rect 499 -561 533 -527
rect 499 -629 533 -595
rect 499 -697 533 -663
rect 499 -765 533 -731
rect 499 -833 533 -799
rect 499 -901 533 -867
rect 499 -969 533 -935
rect 499 -1037 533 -1003
rect 499 -1105 533 -1071
rect 499 -1173 533 -1139
rect 499 -1241 533 -1207
rect 499 -1309 533 -1275
rect 499 -1377 533 -1343
rect 499 -1445 533 -1411
rect 499 -1513 533 -1479
rect 499 -1581 533 -1547
rect 499 -1649 533 -1615
rect 499 -1717 533 -1683
rect 499 -1785 533 -1751
rect 499 -1853 533 -1819
rect 499 -1921 533 -1887
rect 499 -1989 533 -1955
rect 499 -2057 533 -2023
rect 499 -2125 533 -2091
rect 499 -2193 533 -2159
rect 499 -2261 533 -2227
rect 499 -2329 533 -2295
rect 499 -2397 533 -2363
rect 499 -2465 533 -2431
rect 757 2431 791 2465
rect 757 2363 791 2397
rect 757 2295 791 2329
rect 757 2227 791 2261
rect 757 2159 791 2193
rect 757 2091 791 2125
rect 757 2023 791 2057
rect 757 1955 791 1989
rect 757 1887 791 1921
rect 757 1819 791 1853
rect 757 1751 791 1785
rect 757 1683 791 1717
rect 757 1615 791 1649
rect 757 1547 791 1581
rect 757 1479 791 1513
rect 757 1411 791 1445
rect 757 1343 791 1377
rect 757 1275 791 1309
rect 757 1207 791 1241
rect 757 1139 791 1173
rect 757 1071 791 1105
rect 757 1003 791 1037
rect 757 935 791 969
rect 757 867 791 901
rect 757 799 791 833
rect 757 731 791 765
rect 757 663 791 697
rect 757 595 791 629
rect 757 527 791 561
rect 757 459 791 493
rect 757 391 791 425
rect 757 323 791 357
rect 757 255 791 289
rect 757 187 791 221
rect 757 119 791 153
rect 757 51 791 85
rect 757 -17 791 17
rect 757 -85 791 -51
rect 757 -153 791 -119
rect 757 -221 791 -187
rect 757 -289 791 -255
rect 757 -357 791 -323
rect 757 -425 791 -391
rect 757 -493 791 -459
rect 757 -561 791 -527
rect 757 -629 791 -595
rect 757 -697 791 -663
rect 757 -765 791 -731
rect 757 -833 791 -799
rect 757 -901 791 -867
rect 757 -969 791 -935
rect 757 -1037 791 -1003
rect 757 -1105 791 -1071
rect 757 -1173 791 -1139
rect 757 -1241 791 -1207
rect 757 -1309 791 -1275
rect 757 -1377 791 -1343
rect 757 -1445 791 -1411
rect 757 -1513 791 -1479
rect 757 -1581 791 -1547
rect 757 -1649 791 -1615
rect 757 -1717 791 -1683
rect 757 -1785 791 -1751
rect 757 -1853 791 -1819
rect 757 -1921 791 -1887
rect 757 -1989 791 -1955
rect 757 -2057 791 -2023
rect 757 -2125 791 -2091
rect 757 -2193 791 -2159
rect 757 -2261 791 -2227
rect 757 -2329 791 -2295
rect 757 -2397 791 -2363
rect 757 -2465 791 -2431
rect 1015 2431 1049 2465
rect 1015 2363 1049 2397
rect 1015 2295 1049 2329
rect 1015 2227 1049 2261
rect 1015 2159 1049 2193
rect 1015 2091 1049 2125
rect 1015 2023 1049 2057
rect 1015 1955 1049 1989
rect 1015 1887 1049 1921
rect 1015 1819 1049 1853
rect 1015 1751 1049 1785
rect 1015 1683 1049 1717
rect 1015 1615 1049 1649
rect 1015 1547 1049 1581
rect 1015 1479 1049 1513
rect 1015 1411 1049 1445
rect 1015 1343 1049 1377
rect 1015 1275 1049 1309
rect 1015 1207 1049 1241
rect 1015 1139 1049 1173
rect 1015 1071 1049 1105
rect 1015 1003 1049 1037
rect 1015 935 1049 969
rect 1015 867 1049 901
rect 1015 799 1049 833
rect 1015 731 1049 765
rect 1015 663 1049 697
rect 1015 595 1049 629
rect 1015 527 1049 561
rect 1015 459 1049 493
rect 1015 391 1049 425
rect 1015 323 1049 357
rect 1015 255 1049 289
rect 1015 187 1049 221
rect 1015 119 1049 153
rect 1015 51 1049 85
rect 1015 -17 1049 17
rect 1015 -85 1049 -51
rect 1015 -153 1049 -119
rect 1015 -221 1049 -187
rect 1015 -289 1049 -255
rect 1015 -357 1049 -323
rect 1015 -425 1049 -391
rect 1015 -493 1049 -459
rect 1015 -561 1049 -527
rect 1015 -629 1049 -595
rect 1015 -697 1049 -663
rect 1015 -765 1049 -731
rect 1015 -833 1049 -799
rect 1015 -901 1049 -867
rect 1015 -969 1049 -935
rect 1015 -1037 1049 -1003
rect 1015 -1105 1049 -1071
rect 1015 -1173 1049 -1139
rect 1015 -1241 1049 -1207
rect 1015 -1309 1049 -1275
rect 1015 -1377 1049 -1343
rect 1015 -1445 1049 -1411
rect 1015 -1513 1049 -1479
rect 1015 -1581 1049 -1547
rect 1015 -1649 1049 -1615
rect 1015 -1717 1049 -1683
rect 1015 -1785 1049 -1751
rect 1015 -1853 1049 -1819
rect 1015 -1921 1049 -1887
rect 1015 -1989 1049 -1955
rect 1015 -2057 1049 -2023
rect 1015 -2125 1049 -2091
rect 1015 -2193 1049 -2159
rect 1015 -2261 1049 -2227
rect 1015 -2329 1049 -2295
rect 1015 -2397 1049 -2363
rect 1015 -2465 1049 -2431
rect 1273 2431 1307 2465
rect 1273 2363 1307 2397
rect 1273 2295 1307 2329
rect 1273 2227 1307 2261
rect 1273 2159 1307 2193
rect 1273 2091 1307 2125
rect 1273 2023 1307 2057
rect 1273 1955 1307 1989
rect 1273 1887 1307 1921
rect 1273 1819 1307 1853
rect 1273 1751 1307 1785
rect 1273 1683 1307 1717
rect 1273 1615 1307 1649
rect 1273 1547 1307 1581
rect 1273 1479 1307 1513
rect 1273 1411 1307 1445
rect 1273 1343 1307 1377
rect 1273 1275 1307 1309
rect 1273 1207 1307 1241
rect 1273 1139 1307 1173
rect 1273 1071 1307 1105
rect 1273 1003 1307 1037
rect 1273 935 1307 969
rect 1273 867 1307 901
rect 1273 799 1307 833
rect 1273 731 1307 765
rect 1273 663 1307 697
rect 1273 595 1307 629
rect 1273 527 1307 561
rect 1273 459 1307 493
rect 1273 391 1307 425
rect 1273 323 1307 357
rect 1273 255 1307 289
rect 1273 187 1307 221
rect 1273 119 1307 153
rect 1273 51 1307 85
rect 1273 -17 1307 17
rect 1273 -85 1307 -51
rect 1273 -153 1307 -119
rect 1273 -221 1307 -187
rect 1273 -289 1307 -255
rect 1273 -357 1307 -323
rect 1273 -425 1307 -391
rect 1273 -493 1307 -459
rect 1273 -561 1307 -527
rect 1273 -629 1307 -595
rect 1273 -697 1307 -663
rect 1273 -765 1307 -731
rect 1273 -833 1307 -799
rect 1273 -901 1307 -867
rect 1273 -969 1307 -935
rect 1273 -1037 1307 -1003
rect 1273 -1105 1307 -1071
rect 1273 -1173 1307 -1139
rect 1273 -1241 1307 -1207
rect 1273 -1309 1307 -1275
rect 1273 -1377 1307 -1343
rect 1273 -1445 1307 -1411
rect 1273 -1513 1307 -1479
rect 1273 -1581 1307 -1547
rect 1273 -1649 1307 -1615
rect 1273 -1717 1307 -1683
rect 1273 -1785 1307 -1751
rect 1273 -1853 1307 -1819
rect 1273 -1921 1307 -1887
rect 1273 -1989 1307 -1955
rect 1273 -2057 1307 -2023
rect 1273 -2125 1307 -2091
rect 1273 -2193 1307 -2159
rect 1273 -2261 1307 -2227
rect 1273 -2329 1307 -2295
rect 1273 -2397 1307 -2363
rect 1273 -2465 1307 -2431
<< psubdiff >>
rect -1421 2640 -1309 2674
rect -1275 2640 -1241 2674
rect -1207 2640 -1173 2674
rect -1139 2640 -1105 2674
rect -1071 2640 -1037 2674
rect -1003 2640 -969 2674
rect -935 2640 -901 2674
rect -867 2640 -833 2674
rect -799 2640 -765 2674
rect -731 2640 -697 2674
rect -663 2640 -629 2674
rect -595 2640 -561 2674
rect -527 2640 -493 2674
rect -459 2640 -425 2674
rect -391 2640 -357 2674
rect -323 2640 -289 2674
rect -255 2640 -221 2674
rect -187 2640 -153 2674
rect -119 2640 -85 2674
rect -51 2640 -17 2674
rect 17 2640 51 2674
rect 85 2640 119 2674
rect 153 2640 187 2674
rect 221 2640 255 2674
rect 289 2640 323 2674
rect 357 2640 391 2674
rect 425 2640 459 2674
rect 493 2640 527 2674
rect 561 2640 595 2674
rect 629 2640 663 2674
rect 697 2640 731 2674
rect 765 2640 799 2674
rect 833 2640 867 2674
rect 901 2640 935 2674
rect 969 2640 1003 2674
rect 1037 2640 1071 2674
rect 1105 2640 1139 2674
rect 1173 2640 1207 2674
rect 1241 2640 1275 2674
rect 1309 2640 1421 2674
rect -1421 2567 -1387 2640
rect -1421 2499 -1387 2533
rect 1387 2567 1421 2640
rect -1421 2431 -1387 2465
rect -1421 2363 -1387 2397
rect -1421 2295 -1387 2329
rect -1421 2227 -1387 2261
rect -1421 2159 -1387 2193
rect -1421 2091 -1387 2125
rect -1421 2023 -1387 2057
rect -1421 1955 -1387 1989
rect -1421 1887 -1387 1921
rect -1421 1819 -1387 1853
rect -1421 1751 -1387 1785
rect -1421 1683 -1387 1717
rect -1421 1615 -1387 1649
rect -1421 1547 -1387 1581
rect -1421 1479 -1387 1513
rect -1421 1411 -1387 1445
rect -1421 1343 -1387 1377
rect -1421 1275 -1387 1309
rect -1421 1207 -1387 1241
rect -1421 1139 -1387 1173
rect -1421 1071 -1387 1105
rect -1421 1003 -1387 1037
rect -1421 935 -1387 969
rect -1421 867 -1387 901
rect -1421 799 -1387 833
rect -1421 731 -1387 765
rect -1421 663 -1387 697
rect -1421 595 -1387 629
rect -1421 527 -1387 561
rect -1421 459 -1387 493
rect -1421 391 -1387 425
rect -1421 323 -1387 357
rect -1421 255 -1387 289
rect -1421 187 -1387 221
rect -1421 119 -1387 153
rect -1421 51 -1387 85
rect -1421 -17 -1387 17
rect -1421 -85 -1387 -51
rect -1421 -153 -1387 -119
rect -1421 -221 -1387 -187
rect -1421 -289 -1387 -255
rect -1421 -357 -1387 -323
rect -1421 -425 -1387 -391
rect -1421 -493 -1387 -459
rect -1421 -561 -1387 -527
rect -1421 -629 -1387 -595
rect -1421 -697 -1387 -663
rect -1421 -765 -1387 -731
rect -1421 -833 -1387 -799
rect -1421 -901 -1387 -867
rect -1421 -969 -1387 -935
rect -1421 -1037 -1387 -1003
rect -1421 -1105 -1387 -1071
rect -1421 -1173 -1387 -1139
rect -1421 -1241 -1387 -1207
rect -1421 -1309 -1387 -1275
rect -1421 -1377 -1387 -1343
rect -1421 -1445 -1387 -1411
rect -1421 -1513 -1387 -1479
rect -1421 -1581 -1387 -1547
rect -1421 -1649 -1387 -1615
rect -1421 -1717 -1387 -1683
rect -1421 -1785 -1387 -1751
rect -1421 -1853 -1387 -1819
rect -1421 -1921 -1387 -1887
rect -1421 -1989 -1387 -1955
rect -1421 -2057 -1387 -2023
rect -1421 -2125 -1387 -2091
rect -1421 -2193 -1387 -2159
rect -1421 -2261 -1387 -2227
rect -1421 -2329 -1387 -2295
rect -1421 -2397 -1387 -2363
rect -1421 -2465 -1387 -2431
rect -1421 -2533 -1387 -2499
rect 1387 2499 1421 2533
rect 1387 2431 1421 2465
rect 1387 2363 1421 2397
rect 1387 2295 1421 2329
rect 1387 2227 1421 2261
rect 1387 2159 1421 2193
rect 1387 2091 1421 2125
rect 1387 2023 1421 2057
rect 1387 1955 1421 1989
rect 1387 1887 1421 1921
rect 1387 1819 1421 1853
rect 1387 1751 1421 1785
rect 1387 1683 1421 1717
rect 1387 1615 1421 1649
rect 1387 1547 1421 1581
rect 1387 1479 1421 1513
rect 1387 1411 1421 1445
rect 1387 1343 1421 1377
rect 1387 1275 1421 1309
rect 1387 1207 1421 1241
rect 1387 1139 1421 1173
rect 1387 1071 1421 1105
rect 1387 1003 1421 1037
rect 1387 935 1421 969
rect 1387 867 1421 901
rect 1387 799 1421 833
rect 1387 731 1421 765
rect 1387 663 1421 697
rect 1387 595 1421 629
rect 1387 527 1421 561
rect 1387 459 1421 493
rect 1387 391 1421 425
rect 1387 323 1421 357
rect 1387 255 1421 289
rect 1387 187 1421 221
rect 1387 119 1421 153
rect 1387 51 1421 85
rect 1387 -17 1421 17
rect 1387 -85 1421 -51
rect 1387 -153 1421 -119
rect 1387 -221 1421 -187
rect 1387 -289 1421 -255
rect 1387 -357 1421 -323
rect 1387 -425 1421 -391
rect 1387 -493 1421 -459
rect 1387 -561 1421 -527
rect 1387 -629 1421 -595
rect 1387 -697 1421 -663
rect 1387 -765 1421 -731
rect 1387 -833 1421 -799
rect 1387 -901 1421 -867
rect 1387 -969 1421 -935
rect 1387 -1037 1421 -1003
rect 1387 -1105 1421 -1071
rect 1387 -1173 1421 -1139
rect 1387 -1241 1421 -1207
rect 1387 -1309 1421 -1275
rect 1387 -1377 1421 -1343
rect 1387 -1445 1421 -1411
rect 1387 -1513 1421 -1479
rect 1387 -1581 1421 -1547
rect 1387 -1649 1421 -1615
rect 1387 -1717 1421 -1683
rect 1387 -1785 1421 -1751
rect 1387 -1853 1421 -1819
rect 1387 -1921 1421 -1887
rect 1387 -1989 1421 -1955
rect 1387 -2057 1421 -2023
rect 1387 -2125 1421 -2091
rect 1387 -2193 1421 -2159
rect 1387 -2261 1421 -2227
rect 1387 -2329 1421 -2295
rect 1387 -2397 1421 -2363
rect 1387 -2465 1421 -2431
rect -1421 -2640 -1387 -2567
rect 1387 -2533 1421 -2499
rect 1387 -2640 1421 -2567
rect -1421 -2674 -1309 -2640
rect -1275 -2674 -1241 -2640
rect -1207 -2674 -1173 -2640
rect -1139 -2674 -1105 -2640
rect -1071 -2674 -1037 -2640
rect -1003 -2674 -969 -2640
rect -935 -2674 -901 -2640
rect -867 -2674 -833 -2640
rect -799 -2674 -765 -2640
rect -731 -2674 -697 -2640
rect -663 -2674 -629 -2640
rect -595 -2674 -561 -2640
rect -527 -2674 -493 -2640
rect -459 -2674 -425 -2640
rect -391 -2674 -357 -2640
rect -323 -2674 -289 -2640
rect -255 -2674 -221 -2640
rect -187 -2674 -153 -2640
rect -119 -2674 -85 -2640
rect -51 -2674 -17 -2640
rect 17 -2674 51 -2640
rect 85 -2674 119 -2640
rect 153 -2674 187 -2640
rect 221 -2674 255 -2640
rect 289 -2674 323 -2640
rect 357 -2674 391 -2640
rect 425 -2674 459 -2640
rect 493 -2674 527 -2640
rect 561 -2674 595 -2640
rect 629 -2674 663 -2640
rect 697 -2674 731 -2640
rect 765 -2674 799 -2640
rect 833 -2674 867 -2640
rect 901 -2674 935 -2640
rect 969 -2674 1003 -2640
rect 1037 -2674 1071 -2640
rect 1105 -2674 1139 -2640
rect 1173 -2674 1207 -2640
rect 1241 -2674 1275 -2640
rect 1309 -2674 1421 -2640
<< psubdiffcont >>
rect -1309 2640 -1275 2674
rect -1241 2640 -1207 2674
rect -1173 2640 -1139 2674
rect -1105 2640 -1071 2674
rect -1037 2640 -1003 2674
rect -969 2640 -935 2674
rect -901 2640 -867 2674
rect -833 2640 -799 2674
rect -765 2640 -731 2674
rect -697 2640 -663 2674
rect -629 2640 -595 2674
rect -561 2640 -527 2674
rect -493 2640 -459 2674
rect -425 2640 -391 2674
rect -357 2640 -323 2674
rect -289 2640 -255 2674
rect -221 2640 -187 2674
rect -153 2640 -119 2674
rect -85 2640 -51 2674
rect -17 2640 17 2674
rect 51 2640 85 2674
rect 119 2640 153 2674
rect 187 2640 221 2674
rect 255 2640 289 2674
rect 323 2640 357 2674
rect 391 2640 425 2674
rect 459 2640 493 2674
rect 527 2640 561 2674
rect 595 2640 629 2674
rect 663 2640 697 2674
rect 731 2640 765 2674
rect 799 2640 833 2674
rect 867 2640 901 2674
rect 935 2640 969 2674
rect 1003 2640 1037 2674
rect 1071 2640 1105 2674
rect 1139 2640 1173 2674
rect 1207 2640 1241 2674
rect 1275 2640 1309 2674
rect -1421 2533 -1387 2567
rect 1387 2533 1421 2567
rect -1421 2465 -1387 2499
rect -1421 2397 -1387 2431
rect -1421 2329 -1387 2363
rect -1421 2261 -1387 2295
rect -1421 2193 -1387 2227
rect -1421 2125 -1387 2159
rect -1421 2057 -1387 2091
rect -1421 1989 -1387 2023
rect -1421 1921 -1387 1955
rect -1421 1853 -1387 1887
rect -1421 1785 -1387 1819
rect -1421 1717 -1387 1751
rect -1421 1649 -1387 1683
rect -1421 1581 -1387 1615
rect -1421 1513 -1387 1547
rect -1421 1445 -1387 1479
rect -1421 1377 -1387 1411
rect -1421 1309 -1387 1343
rect -1421 1241 -1387 1275
rect -1421 1173 -1387 1207
rect -1421 1105 -1387 1139
rect -1421 1037 -1387 1071
rect -1421 969 -1387 1003
rect -1421 901 -1387 935
rect -1421 833 -1387 867
rect -1421 765 -1387 799
rect -1421 697 -1387 731
rect -1421 629 -1387 663
rect -1421 561 -1387 595
rect -1421 493 -1387 527
rect -1421 425 -1387 459
rect -1421 357 -1387 391
rect -1421 289 -1387 323
rect -1421 221 -1387 255
rect -1421 153 -1387 187
rect -1421 85 -1387 119
rect -1421 17 -1387 51
rect -1421 -51 -1387 -17
rect -1421 -119 -1387 -85
rect -1421 -187 -1387 -153
rect -1421 -255 -1387 -221
rect -1421 -323 -1387 -289
rect -1421 -391 -1387 -357
rect -1421 -459 -1387 -425
rect -1421 -527 -1387 -493
rect -1421 -595 -1387 -561
rect -1421 -663 -1387 -629
rect -1421 -731 -1387 -697
rect -1421 -799 -1387 -765
rect -1421 -867 -1387 -833
rect -1421 -935 -1387 -901
rect -1421 -1003 -1387 -969
rect -1421 -1071 -1387 -1037
rect -1421 -1139 -1387 -1105
rect -1421 -1207 -1387 -1173
rect -1421 -1275 -1387 -1241
rect -1421 -1343 -1387 -1309
rect -1421 -1411 -1387 -1377
rect -1421 -1479 -1387 -1445
rect -1421 -1547 -1387 -1513
rect -1421 -1615 -1387 -1581
rect -1421 -1683 -1387 -1649
rect -1421 -1751 -1387 -1717
rect -1421 -1819 -1387 -1785
rect -1421 -1887 -1387 -1853
rect -1421 -1955 -1387 -1921
rect -1421 -2023 -1387 -1989
rect -1421 -2091 -1387 -2057
rect -1421 -2159 -1387 -2125
rect -1421 -2227 -1387 -2193
rect -1421 -2295 -1387 -2261
rect -1421 -2363 -1387 -2329
rect -1421 -2431 -1387 -2397
rect -1421 -2499 -1387 -2465
rect 1387 2465 1421 2499
rect 1387 2397 1421 2431
rect 1387 2329 1421 2363
rect 1387 2261 1421 2295
rect 1387 2193 1421 2227
rect 1387 2125 1421 2159
rect 1387 2057 1421 2091
rect 1387 1989 1421 2023
rect 1387 1921 1421 1955
rect 1387 1853 1421 1887
rect 1387 1785 1421 1819
rect 1387 1717 1421 1751
rect 1387 1649 1421 1683
rect 1387 1581 1421 1615
rect 1387 1513 1421 1547
rect 1387 1445 1421 1479
rect 1387 1377 1421 1411
rect 1387 1309 1421 1343
rect 1387 1241 1421 1275
rect 1387 1173 1421 1207
rect 1387 1105 1421 1139
rect 1387 1037 1421 1071
rect 1387 969 1421 1003
rect 1387 901 1421 935
rect 1387 833 1421 867
rect 1387 765 1421 799
rect 1387 697 1421 731
rect 1387 629 1421 663
rect 1387 561 1421 595
rect 1387 493 1421 527
rect 1387 425 1421 459
rect 1387 357 1421 391
rect 1387 289 1421 323
rect 1387 221 1421 255
rect 1387 153 1421 187
rect 1387 85 1421 119
rect 1387 17 1421 51
rect 1387 -51 1421 -17
rect 1387 -119 1421 -85
rect 1387 -187 1421 -153
rect 1387 -255 1421 -221
rect 1387 -323 1421 -289
rect 1387 -391 1421 -357
rect 1387 -459 1421 -425
rect 1387 -527 1421 -493
rect 1387 -595 1421 -561
rect 1387 -663 1421 -629
rect 1387 -731 1421 -697
rect 1387 -799 1421 -765
rect 1387 -867 1421 -833
rect 1387 -935 1421 -901
rect 1387 -1003 1421 -969
rect 1387 -1071 1421 -1037
rect 1387 -1139 1421 -1105
rect 1387 -1207 1421 -1173
rect 1387 -1275 1421 -1241
rect 1387 -1343 1421 -1309
rect 1387 -1411 1421 -1377
rect 1387 -1479 1421 -1445
rect 1387 -1547 1421 -1513
rect 1387 -1615 1421 -1581
rect 1387 -1683 1421 -1649
rect 1387 -1751 1421 -1717
rect 1387 -1819 1421 -1785
rect 1387 -1887 1421 -1853
rect 1387 -1955 1421 -1921
rect 1387 -2023 1421 -1989
rect 1387 -2091 1421 -2057
rect 1387 -2159 1421 -2125
rect 1387 -2227 1421 -2193
rect 1387 -2295 1421 -2261
rect 1387 -2363 1421 -2329
rect 1387 -2431 1421 -2397
rect 1387 -2499 1421 -2465
rect -1421 -2567 -1387 -2533
rect 1387 -2567 1421 -2533
rect -1309 -2674 -1275 -2640
rect -1241 -2674 -1207 -2640
rect -1173 -2674 -1139 -2640
rect -1105 -2674 -1071 -2640
rect -1037 -2674 -1003 -2640
rect -969 -2674 -935 -2640
rect -901 -2674 -867 -2640
rect -833 -2674 -799 -2640
rect -765 -2674 -731 -2640
rect -697 -2674 -663 -2640
rect -629 -2674 -595 -2640
rect -561 -2674 -527 -2640
rect -493 -2674 -459 -2640
rect -425 -2674 -391 -2640
rect -357 -2674 -323 -2640
rect -289 -2674 -255 -2640
rect -221 -2674 -187 -2640
rect -153 -2674 -119 -2640
rect -85 -2674 -51 -2640
rect -17 -2674 17 -2640
rect 51 -2674 85 -2640
rect 119 -2674 153 -2640
rect 187 -2674 221 -2640
rect 255 -2674 289 -2640
rect 323 -2674 357 -2640
rect 391 -2674 425 -2640
rect 459 -2674 493 -2640
rect 527 -2674 561 -2640
rect 595 -2674 629 -2640
rect 663 -2674 697 -2640
rect 731 -2674 765 -2640
rect 799 -2674 833 -2640
rect 867 -2674 901 -2640
rect 935 -2674 969 -2640
rect 1003 -2674 1037 -2640
rect 1071 -2674 1105 -2640
rect 1139 -2674 1173 -2640
rect 1207 -2674 1241 -2640
rect 1275 -2674 1309 -2640
<< poly >>
rect -1261 2572 -1061 2588
rect -1261 2538 -1212 2572
rect -1178 2538 -1144 2572
rect -1110 2538 -1061 2572
rect -1261 2500 -1061 2538
rect -1003 2572 -803 2588
rect -1003 2538 -954 2572
rect -920 2538 -886 2572
rect -852 2538 -803 2572
rect -1003 2500 -803 2538
rect -745 2572 -545 2588
rect -745 2538 -696 2572
rect -662 2538 -628 2572
rect -594 2538 -545 2572
rect -745 2500 -545 2538
rect -487 2572 -287 2588
rect -487 2538 -438 2572
rect -404 2538 -370 2572
rect -336 2538 -287 2572
rect -487 2500 -287 2538
rect -229 2572 -29 2588
rect -229 2538 -180 2572
rect -146 2538 -112 2572
rect -78 2538 -29 2572
rect -229 2500 -29 2538
rect 29 2572 229 2588
rect 29 2538 78 2572
rect 112 2538 146 2572
rect 180 2538 229 2572
rect 29 2500 229 2538
rect 287 2572 487 2588
rect 287 2538 336 2572
rect 370 2538 404 2572
rect 438 2538 487 2572
rect 287 2500 487 2538
rect 545 2572 745 2588
rect 545 2538 594 2572
rect 628 2538 662 2572
rect 696 2538 745 2572
rect 545 2500 745 2538
rect 803 2572 1003 2588
rect 803 2538 852 2572
rect 886 2538 920 2572
rect 954 2538 1003 2572
rect 803 2500 1003 2538
rect 1061 2572 1261 2588
rect 1061 2538 1110 2572
rect 1144 2538 1178 2572
rect 1212 2538 1261 2572
rect 1061 2500 1261 2538
rect -1261 -2538 -1061 -2500
rect -1261 -2572 -1212 -2538
rect -1178 -2572 -1144 -2538
rect -1110 -2572 -1061 -2538
rect -1261 -2588 -1061 -2572
rect -1003 -2538 -803 -2500
rect -1003 -2572 -954 -2538
rect -920 -2572 -886 -2538
rect -852 -2572 -803 -2538
rect -1003 -2588 -803 -2572
rect -745 -2538 -545 -2500
rect -745 -2572 -696 -2538
rect -662 -2572 -628 -2538
rect -594 -2572 -545 -2538
rect -745 -2588 -545 -2572
rect -487 -2538 -287 -2500
rect -487 -2572 -438 -2538
rect -404 -2572 -370 -2538
rect -336 -2572 -287 -2538
rect -487 -2588 -287 -2572
rect -229 -2538 -29 -2500
rect -229 -2572 -180 -2538
rect -146 -2572 -112 -2538
rect -78 -2572 -29 -2538
rect -229 -2588 -29 -2572
rect 29 -2538 229 -2500
rect 29 -2572 78 -2538
rect 112 -2572 146 -2538
rect 180 -2572 229 -2538
rect 29 -2588 229 -2572
rect 287 -2538 487 -2500
rect 287 -2572 336 -2538
rect 370 -2572 404 -2538
rect 438 -2572 487 -2538
rect 287 -2588 487 -2572
rect 545 -2538 745 -2500
rect 545 -2572 594 -2538
rect 628 -2572 662 -2538
rect 696 -2572 745 -2538
rect 545 -2588 745 -2572
rect 803 -2538 1003 -2500
rect 803 -2572 852 -2538
rect 886 -2572 920 -2538
rect 954 -2572 1003 -2538
rect 803 -2588 1003 -2572
rect 1061 -2538 1261 -2500
rect 1061 -2572 1110 -2538
rect 1144 -2572 1178 -2538
rect 1212 -2572 1261 -2538
rect 1061 -2588 1261 -2572
<< polycont >>
rect -1212 2538 -1178 2572
rect -1144 2538 -1110 2572
rect -954 2538 -920 2572
rect -886 2538 -852 2572
rect -696 2538 -662 2572
rect -628 2538 -594 2572
rect -438 2538 -404 2572
rect -370 2538 -336 2572
rect -180 2538 -146 2572
rect -112 2538 -78 2572
rect 78 2538 112 2572
rect 146 2538 180 2572
rect 336 2538 370 2572
rect 404 2538 438 2572
rect 594 2538 628 2572
rect 662 2538 696 2572
rect 852 2538 886 2572
rect 920 2538 954 2572
rect 1110 2538 1144 2572
rect 1178 2538 1212 2572
rect -1212 -2572 -1178 -2538
rect -1144 -2572 -1110 -2538
rect -954 -2572 -920 -2538
rect -886 -2572 -852 -2538
rect -696 -2572 -662 -2538
rect -628 -2572 -594 -2538
rect -438 -2572 -404 -2538
rect -370 -2572 -336 -2538
rect -180 -2572 -146 -2538
rect -112 -2572 -78 -2538
rect 78 -2572 112 -2538
rect 146 -2572 180 -2538
rect 336 -2572 370 -2538
rect 404 -2572 438 -2538
rect 594 -2572 628 -2538
rect 662 -2572 696 -2538
rect 852 -2572 886 -2538
rect 920 -2572 954 -2538
rect 1110 -2572 1144 -2538
rect 1178 -2572 1212 -2538
<< locali >>
rect -1421 2640 -1309 2674
rect -1275 2640 -1241 2674
rect -1207 2640 -1173 2674
rect -1139 2640 -1105 2674
rect -1071 2640 -1037 2674
rect -1003 2640 -969 2674
rect -935 2640 -901 2674
rect -867 2640 -833 2674
rect -799 2640 -765 2674
rect -731 2640 -697 2674
rect -663 2640 -629 2674
rect -595 2640 -561 2674
rect -527 2640 -493 2674
rect -459 2640 -425 2674
rect -391 2640 -357 2674
rect -323 2640 -289 2674
rect -255 2640 -221 2674
rect -187 2640 -153 2674
rect -119 2640 -85 2674
rect -51 2640 -17 2674
rect 17 2640 51 2674
rect 85 2640 119 2674
rect 153 2640 187 2674
rect 221 2640 255 2674
rect 289 2640 323 2674
rect 357 2640 391 2674
rect 425 2640 459 2674
rect 493 2640 527 2674
rect 561 2640 595 2674
rect 629 2640 663 2674
rect 697 2640 731 2674
rect 765 2640 799 2674
rect 833 2640 867 2674
rect 901 2640 935 2674
rect 969 2640 1003 2674
rect 1037 2640 1071 2674
rect 1105 2640 1139 2674
rect 1173 2640 1207 2674
rect 1241 2640 1275 2674
rect 1309 2640 1421 2674
rect -1421 2567 -1387 2640
rect -1261 2538 -1214 2572
rect -1178 2538 -1144 2572
rect -1108 2538 -1061 2572
rect -1003 2538 -956 2572
rect -920 2538 -886 2572
rect -850 2538 -803 2572
rect -745 2538 -698 2572
rect -662 2538 -628 2572
rect -592 2538 -545 2572
rect -487 2538 -440 2572
rect -404 2538 -370 2572
rect -334 2538 -287 2572
rect -229 2538 -182 2572
rect -146 2538 -112 2572
rect -76 2538 -29 2572
rect 29 2538 76 2572
rect 112 2538 146 2572
rect 182 2538 229 2572
rect 287 2538 334 2572
rect 370 2538 404 2572
rect 440 2538 487 2572
rect 545 2538 592 2572
rect 628 2538 662 2572
rect 698 2538 745 2572
rect 803 2538 850 2572
rect 886 2538 920 2572
rect 956 2538 1003 2572
rect 1061 2538 1108 2572
rect 1144 2538 1178 2572
rect 1214 2538 1261 2572
rect 1387 2567 1421 2640
rect -1421 2499 -1387 2533
rect -1421 2431 -1387 2465
rect -1421 2363 -1387 2397
rect -1421 2295 -1387 2329
rect -1421 2227 -1387 2261
rect -1421 2159 -1387 2193
rect -1421 2091 -1387 2125
rect -1421 2023 -1387 2057
rect -1421 1955 -1387 1989
rect -1421 1887 -1387 1921
rect -1421 1819 -1387 1853
rect -1421 1751 -1387 1785
rect -1421 1683 -1387 1717
rect -1421 1615 -1387 1649
rect -1421 1547 -1387 1581
rect -1421 1479 -1387 1513
rect -1421 1411 -1387 1445
rect -1421 1343 -1387 1377
rect -1421 1275 -1387 1309
rect -1421 1207 -1387 1241
rect -1421 1139 -1387 1173
rect -1421 1071 -1387 1105
rect -1421 1003 -1387 1037
rect -1421 935 -1387 969
rect -1421 867 -1387 901
rect -1421 799 -1387 833
rect -1421 731 -1387 765
rect -1421 663 -1387 697
rect -1421 595 -1387 629
rect -1421 527 -1387 561
rect -1421 459 -1387 493
rect -1421 391 -1387 425
rect -1421 323 -1387 357
rect -1421 255 -1387 289
rect -1421 187 -1387 221
rect -1421 119 -1387 153
rect -1421 51 -1387 85
rect -1421 -17 -1387 17
rect -1421 -85 -1387 -51
rect -1421 -153 -1387 -119
rect -1421 -221 -1387 -187
rect -1421 -289 -1387 -255
rect -1421 -357 -1387 -323
rect -1421 -425 -1387 -391
rect -1421 -493 -1387 -459
rect -1421 -561 -1387 -527
rect -1421 -629 -1387 -595
rect -1421 -697 -1387 -663
rect -1421 -765 -1387 -731
rect -1421 -833 -1387 -799
rect -1421 -901 -1387 -867
rect -1421 -969 -1387 -935
rect -1421 -1037 -1387 -1003
rect -1421 -1105 -1387 -1071
rect -1421 -1173 -1387 -1139
rect -1421 -1241 -1387 -1207
rect -1421 -1309 -1387 -1275
rect -1421 -1377 -1387 -1343
rect -1421 -1445 -1387 -1411
rect -1421 -1513 -1387 -1479
rect -1421 -1581 -1387 -1547
rect -1421 -1649 -1387 -1615
rect -1421 -1717 -1387 -1683
rect -1421 -1785 -1387 -1751
rect -1421 -1853 -1387 -1819
rect -1421 -1921 -1387 -1887
rect -1421 -1989 -1387 -1955
rect -1421 -2057 -1387 -2023
rect -1421 -2125 -1387 -2091
rect -1421 -2193 -1387 -2159
rect -1421 -2261 -1387 -2227
rect -1421 -2329 -1387 -2295
rect -1421 -2397 -1387 -2363
rect -1421 -2465 -1387 -2431
rect -1421 -2533 -1387 -2499
rect -1307 2465 -1273 2504
rect -1307 2397 -1273 2431
rect -1307 2329 -1273 2359
rect -1307 2261 -1273 2287
rect -1307 2193 -1273 2215
rect -1307 2125 -1273 2143
rect -1307 2057 -1273 2071
rect -1307 1989 -1273 1999
rect -1307 1921 -1273 1927
rect -1307 1853 -1273 1855
rect -1307 1817 -1273 1819
rect -1307 1745 -1273 1751
rect -1307 1673 -1273 1683
rect -1307 1601 -1273 1615
rect -1307 1529 -1273 1547
rect -1307 1457 -1273 1479
rect -1307 1385 -1273 1411
rect -1307 1313 -1273 1343
rect -1307 1241 -1273 1275
rect -1307 1173 -1273 1207
rect -1307 1105 -1273 1135
rect -1307 1037 -1273 1063
rect -1307 969 -1273 991
rect -1307 901 -1273 919
rect -1307 833 -1273 847
rect -1307 765 -1273 775
rect -1307 697 -1273 703
rect -1307 629 -1273 631
rect -1307 593 -1273 595
rect -1307 521 -1273 527
rect -1307 449 -1273 459
rect -1307 377 -1273 391
rect -1307 305 -1273 323
rect -1307 233 -1273 255
rect -1307 161 -1273 187
rect -1307 89 -1273 119
rect -1307 17 -1273 51
rect -1307 -51 -1273 -17
rect -1307 -119 -1273 -89
rect -1307 -187 -1273 -161
rect -1307 -255 -1273 -233
rect -1307 -323 -1273 -305
rect -1307 -391 -1273 -377
rect -1307 -459 -1273 -449
rect -1307 -527 -1273 -521
rect -1307 -595 -1273 -593
rect -1307 -631 -1273 -629
rect -1307 -703 -1273 -697
rect -1307 -775 -1273 -765
rect -1307 -847 -1273 -833
rect -1307 -919 -1273 -901
rect -1307 -991 -1273 -969
rect -1307 -1063 -1273 -1037
rect -1307 -1135 -1273 -1105
rect -1307 -1207 -1273 -1173
rect -1307 -1275 -1273 -1241
rect -1307 -1343 -1273 -1313
rect -1307 -1411 -1273 -1385
rect -1307 -1479 -1273 -1457
rect -1307 -1547 -1273 -1529
rect -1307 -1615 -1273 -1601
rect -1307 -1683 -1273 -1673
rect -1307 -1751 -1273 -1745
rect -1307 -1819 -1273 -1817
rect -1307 -1855 -1273 -1853
rect -1307 -1927 -1273 -1921
rect -1307 -1999 -1273 -1989
rect -1307 -2071 -1273 -2057
rect -1307 -2143 -1273 -2125
rect -1307 -2215 -1273 -2193
rect -1307 -2287 -1273 -2261
rect -1307 -2359 -1273 -2329
rect -1307 -2431 -1273 -2397
rect -1307 -2504 -1273 -2465
rect -1049 2465 -1015 2504
rect -1049 2397 -1015 2431
rect -1049 2329 -1015 2359
rect -1049 2261 -1015 2287
rect -1049 2193 -1015 2215
rect -1049 2125 -1015 2143
rect -1049 2057 -1015 2071
rect -1049 1989 -1015 1999
rect -1049 1921 -1015 1927
rect -1049 1853 -1015 1855
rect -1049 1817 -1015 1819
rect -1049 1745 -1015 1751
rect -1049 1673 -1015 1683
rect -1049 1601 -1015 1615
rect -1049 1529 -1015 1547
rect -1049 1457 -1015 1479
rect -1049 1385 -1015 1411
rect -1049 1313 -1015 1343
rect -1049 1241 -1015 1275
rect -1049 1173 -1015 1207
rect -1049 1105 -1015 1135
rect -1049 1037 -1015 1063
rect -1049 969 -1015 991
rect -1049 901 -1015 919
rect -1049 833 -1015 847
rect -1049 765 -1015 775
rect -1049 697 -1015 703
rect -1049 629 -1015 631
rect -1049 593 -1015 595
rect -1049 521 -1015 527
rect -1049 449 -1015 459
rect -1049 377 -1015 391
rect -1049 305 -1015 323
rect -1049 233 -1015 255
rect -1049 161 -1015 187
rect -1049 89 -1015 119
rect -1049 17 -1015 51
rect -1049 -51 -1015 -17
rect -1049 -119 -1015 -89
rect -1049 -187 -1015 -161
rect -1049 -255 -1015 -233
rect -1049 -323 -1015 -305
rect -1049 -391 -1015 -377
rect -1049 -459 -1015 -449
rect -1049 -527 -1015 -521
rect -1049 -595 -1015 -593
rect -1049 -631 -1015 -629
rect -1049 -703 -1015 -697
rect -1049 -775 -1015 -765
rect -1049 -847 -1015 -833
rect -1049 -919 -1015 -901
rect -1049 -991 -1015 -969
rect -1049 -1063 -1015 -1037
rect -1049 -1135 -1015 -1105
rect -1049 -1207 -1015 -1173
rect -1049 -1275 -1015 -1241
rect -1049 -1343 -1015 -1313
rect -1049 -1411 -1015 -1385
rect -1049 -1479 -1015 -1457
rect -1049 -1547 -1015 -1529
rect -1049 -1615 -1015 -1601
rect -1049 -1683 -1015 -1673
rect -1049 -1751 -1015 -1745
rect -1049 -1819 -1015 -1817
rect -1049 -1855 -1015 -1853
rect -1049 -1927 -1015 -1921
rect -1049 -1999 -1015 -1989
rect -1049 -2071 -1015 -2057
rect -1049 -2143 -1015 -2125
rect -1049 -2215 -1015 -2193
rect -1049 -2287 -1015 -2261
rect -1049 -2359 -1015 -2329
rect -1049 -2431 -1015 -2397
rect -1049 -2504 -1015 -2465
rect -791 2465 -757 2504
rect -791 2397 -757 2431
rect -791 2329 -757 2359
rect -791 2261 -757 2287
rect -791 2193 -757 2215
rect -791 2125 -757 2143
rect -791 2057 -757 2071
rect -791 1989 -757 1999
rect -791 1921 -757 1927
rect -791 1853 -757 1855
rect -791 1817 -757 1819
rect -791 1745 -757 1751
rect -791 1673 -757 1683
rect -791 1601 -757 1615
rect -791 1529 -757 1547
rect -791 1457 -757 1479
rect -791 1385 -757 1411
rect -791 1313 -757 1343
rect -791 1241 -757 1275
rect -791 1173 -757 1207
rect -791 1105 -757 1135
rect -791 1037 -757 1063
rect -791 969 -757 991
rect -791 901 -757 919
rect -791 833 -757 847
rect -791 765 -757 775
rect -791 697 -757 703
rect -791 629 -757 631
rect -791 593 -757 595
rect -791 521 -757 527
rect -791 449 -757 459
rect -791 377 -757 391
rect -791 305 -757 323
rect -791 233 -757 255
rect -791 161 -757 187
rect -791 89 -757 119
rect -791 17 -757 51
rect -791 -51 -757 -17
rect -791 -119 -757 -89
rect -791 -187 -757 -161
rect -791 -255 -757 -233
rect -791 -323 -757 -305
rect -791 -391 -757 -377
rect -791 -459 -757 -449
rect -791 -527 -757 -521
rect -791 -595 -757 -593
rect -791 -631 -757 -629
rect -791 -703 -757 -697
rect -791 -775 -757 -765
rect -791 -847 -757 -833
rect -791 -919 -757 -901
rect -791 -991 -757 -969
rect -791 -1063 -757 -1037
rect -791 -1135 -757 -1105
rect -791 -1207 -757 -1173
rect -791 -1275 -757 -1241
rect -791 -1343 -757 -1313
rect -791 -1411 -757 -1385
rect -791 -1479 -757 -1457
rect -791 -1547 -757 -1529
rect -791 -1615 -757 -1601
rect -791 -1683 -757 -1673
rect -791 -1751 -757 -1745
rect -791 -1819 -757 -1817
rect -791 -1855 -757 -1853
rect -791 -1927 -757 -1921
rect -791 -1999 -757 -1989
rect -791 -2071 -757 -2057
rect -791 -2143 -757 -2125
rect -791 -2215 -757 -2193
rect -791 -2287 -757 -2261
rect -791 -2359 -757 -2329
rect -791 -2431 -757 -2397
rect -791 -2504 -757 -2465
rect -533 2465 -499 2504
rect -533 2397 -499 2431
rect -533 2329 -499 2359
rect -533 2261 -499 2287
rect -533 2193 -499 2215
rect -533 2125 -499 2143
rect -533 2057 -499 2071
rect -533 1989 -499 1999
rect -533 1921 -499 1927
rect -533 1853 -499 1855
rect -533 1817 -499 1819
rect -533 1745 -499 1751
rect -533 1673 -499 1683
rect -533 1601 -499 1615
rect -533 1529 -499 1547
rect -533 1457 -499 1479
rect -533 1385 -499 1411
rect -533 1313 -499 1343
rect -533 1241 -499 1275
rect -533 1173 -499 1207
rect -533 1105 -499 1135
rect -533 1037 -499 1063
rect -533 969 -499 991
rect -533 901 -499 919
rect -533 833 -499 847
rect -533 765 -499 775
rect -533 697 -499 703
rect -533 629 -499 631
rect -533 593 -499 595
rect -533 521 -499 527
rect -533 449 -499 459
rect -533 377 -499 391
rect -533 305 -499 323
rect -533 233 -499 255
rect -533 161 -499 187
rect -533 89 -499 119
rect -533 17 -499 51
rect -533 -51 -499 -17
rect -533 -119 -499 -89
rect -533 -187 -499 -161
rect -533 -255 -499 -233
rect -533 -323 -499 -305
rect -533 -391 -499 -377
rect -533 -459 -499 -449
rect -533 -527 -499 -521
rect -533 -595 -499 -593
rect -533 -631 -499 -629
rect -533 -703 -499 -697
rect -533 -775 -499 -765
rect -533 -847 -499 -833
rect -533 -919 -499 -901
rect -533 -991 -499 -969
rect -533 -1063 -499 -1037
rect -533 -1135 -499 -1105
rect -533 -1207 -499 -1173
rect -533 -1275 -499 -1241
rect -533 -1343 -499 -1313
rect -533 -1411 -499 -1385
rect -533 -1479 -499 -1457
rect -533 -1547 -499 -1529
rect -533 -1615 -499 -1601
rect -533 -1683 -499 -1673
rect -533 -1751 -499 -1745
rect -533 -1819 -499 -1817
rect -533 -1855 -499 -1853
rect -533 -1927 -499 -1921
rect -533 -1999 -499 -1989
rect -533 -2071 -499 -2057
rect -533 -2143 -499 -2125
rect -533 -2215 -499 -2193
rect -533 -2287 -499 -2261
rect -533 -2359 -499 -2329
rect -533 -2431 -499 -2397
rect -533 -2504 -499 -2465
rect -275 2465 -241 2504
rect -275 2397 -241 2431
rect -275 2329 -241 2359
rect -275 2261 -241 2287
rect -275 2193 -241 2215
rect -275 2125 -241 2143
rect -275 2057 -241 2071
rect -275 1989 -241 1999
rect -275 1921 -241 1927
rect -275 1853 -241 1855
rect -275 1817 -241 1819
rect -275 1745 -241 1751
rect -275 1673 -241 1683
rect -275 1601 -241 1615
rect -275 1529 -241 1547
rect -275 1457 -241 1479
rect -275 1385 -241 1411
rect -275 1313 -241 1343
rect -275 1241 -241 1275
rect -275 1173 -241 1207
rect -275 1105 -241 1135
rect -275 1037 -241 1063
rect -275 969 -241 991
rect -275 901 -241 919
rect -275 833 -241 847
rect -275 765 -241 775
rect -275 697 -241 703
rect -275 629 -241 631
rect -275 593 -241 595
rect -275 521 -241 527
rect -275 449 -241 459
rect -275 377 -241 391
rect -275 305 -241 323
rect -275 233 -241 255
rect -275 161 -241 187
rect -275 89 -241 119
rect -275 17 -241 51
rect -275 -51 -241 -17
rect -275 -119 -241 -89
rect -275 -187 -241 -161
rect -275 -255 -241 -233
rect -275 -323 -241 -305
rect -275 -391 -241 -377
rect -275 -459 -241 -449
rect -275 -527 -241 -521
rect -275 -595 -241 -593
rect -275 -631 -241 -629
rect -275 -703 -241 -697
rect -275 -775 -241 -765
rect -275 -847 -241 -833
rect -275 -919 -241 -901
rect -275 -991 -241 -969
rect -275 -1063 -241 -1037
rect -275 -1135 -241 -1105
rect -275 -1207 -241 -1173
rect -275 -1275 -241 -1241
rect -275 -1343 -241 -1313
rect -275 -1411 -241 -1385
rect -275 -1479 -241 -1457
rect -275 -1547 -241 -1529
rect -275 -1615 -241 -1601
rect -275 -1683 -241 -1673
rect -275 -1751 -241 -1745
rect -275 -1819 -241 -1817
rect -275 -1855 -241 -1853
rect -275 -1927 -241 -1921
rect -275 -1999 -241 -1989
rect -275 -2071 -241 -2057
rect -275 -2143 -241 -2125
rect -275 -2215 -241 -2193
rect -275 -2287 -241 -2261
rect -275 -2359 -241 -2329
rect -275 -2431 -241 -2397
rect -275 -2504 -241 -2465
rect -17 2465 17 2504
rect -17 2397 17 2431
rect -17 2329 17 2359
rect -17 2261 17 2287
rect -17 2193 17 2215
rect -17 2125 17 2143
rect -17 2057 17 2071
rect -17 1989 17 1999
rect -17 1921 17 1927
rect -17 1853 17 1855
rect -17 1817 17 1819
rect -17 1745 17 1751
rect -17 1673 17 1683
rect -17 1601 17 1615
rect -17 1529 17 1547
rect -17 1457 17 1479
rect -17 1385 17 1411
rect -17 1313 17 1343
rect -17 1241 17 1275
rect -17 1173 17 1207
rect -17 1105 17 1135
rect -17 1037 17 1063
rect -17 969 17 991
rect -17 901 17 919
rect -17 833 17 847
rect -17 765 17 775
rect -17 697 17 703
rect -17 629 17 631
rect -17 593 17 595
rect -17 521 17 527
rect -17 449 17 459
rect -17 377 17 391
rect -17 305 17 323
rect -17 233 17 255
rect -17 161 17 187
rect -17 89 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -89
rect -17 -187 17 -161
rect -17 -255 17 -233
rect -17 -323 17 -305
rect -17 -391 17 -377
rect -17 -459 17 -449
rect -17 -527 17 -521
rect -17 -595 17 -593
rect -17 -631 17 -629
rect -17 -703 17 -697
rect -17 -775 17 -765
rect -17 -847 17 -833
rect -17 -919 17 -901
rect -17 -991 17 -969
rect -17 -1063 17 -1037
rect -17 -1135 17 -1105
rect -17 -1207 17 -1173
rect -17 -1275 17 -1241
rect -17 -1343 17 -1313
rect -17 -1411 17 -1385
rect -17 -1479 17 -1457
rect -17 -1547 17 -1529
rect -17 -1615 17 -1601
rect -17 -1683 17 -1673
rect -17 -1751 17 -1745
rect -17 -1819 17 -1817
rect -17 -1855 17 -1853
rect -17 -1927 17 -1921
rect -17 -1999 17 -1989
rect -17 -2071 17 -2057
rect -17 -2143 17 -2125
rect -17 -2215 17 -2193
rect -17 -2287 17 -2261
rect -17 -2359 17 -2329
rect -17 -2431 17 -2397
rect -17 -2504 17 -2465
rect 241 2465 275 2504
rect 241 2397 275 2431
rect 241 2329 275 2359
rect 241 2261 275 2287
rect 241 2193 275 2215
rect 241 2125 275 2143
rect 241 2057 275 2071
rect 241 1989 275 1999
rect 241 1921 275 1927
rect 241 1853 275 1855
rect 241 1817 275 1819
rect 241 1745 275 1751
rect 241 1673 275 1683
rect 241 1601 275 1615
rect 241 1529 275 1547
rect 241 1457 275 1479
rect 241 1385 275 1411
rect 241 1313 275 1343
rect 241 1241 275 1275
rect 241 1173 275 1207
rect 241 1105 275 1135
rect 241 1037 275 1063
rect 241 969 275 991
rect 241 901 275 919
rect 241 833 275 847
rect 241 765 275 775
rect 241 697 275 703
rect 241 629 275 631
rect 241 593 275 595
rect 241 521 275 527
rect 241 449 275 459
rect 241 377 275 391
rect 241 305 275 323
rect 241 233 275 255
rect 241 161 275 187
rect 241 89 275 119
rect 241 17 275 51
rect 241 -51 275 -17
rect 241 -119 275 -89
rect 241 -187 275 -161
rect 241 -255 275 -233
rect 241 -323 275 -305
rect 241 -391 275 -377
rect 241 -459 275 -449
rect 241 -527 275 -521
rect 241 -595 275 -593
rect 241 -631 275 -629
rect 241 -703 275 -697
rect 241 -775 275 -765
rect 241 -847 275 -833
rect 241 -919 275 -901
rect 241 -991 275 -969
rect 241 -1063 275 -1037
rect 241 -1135 275 -1105
rect 241 -1207 275 -1173
rect 241 -1275 275 -1241
rect 241 -1343 275 -1313
rect 241 -1411 275 -1385
rect 241 -1479 275 -1457
rect 241 -1547 275 -1529
rect 241 -1615 275 -1601
rect 241 -1683 275 -1673
rect 241 -1751 275 -1745
rect 241 -1819 275 -1817
rect 241 -1855 275 -1853
rect 241 -1927 275 -1921
rect 241 -1999 275 -1989
rect 241 -2071 275 -2057
rect 241 -2143 275 -2125
rect 241 -2215 275 -2193
rect 241 -2287 275 -2261
rect 241 -2359 275 -2329
rect 241 -2431 275 -2397
rect 241 -2504 275 -2465
rect 499 2465 533 2504
rect 499 2397 533 2431
rect 499 2329 533 2359
rect 499 2261 533 2287
rect 499 2193 533 2215
rect 499 2125 533 2143
rect 499 2057 533 2071
rect 499 1989 533 1999
rect 499 1921 533 1927
rect 499 1853 533 1855
rect 499 1817 533 1819
rect 499 1745 533 1751
rect 499 1673 533 1683
rect 499 1601 533 1615
rect 499 1529 533 1547
rect 499 1457 533 1479
rect 499 1385 533 1411
rect 499 1313 533 1343
rect 499 1241 533 1275
rect 499 1173 533 1207
rect 499 1105 533 1135
rect 499 1037 533 1063
rect 499 969 533 991
rect 499 901 533 919
rect 499 833 533 847
rect 499 765 533 775
rect 499 697 533 703
rect 499 629 533 631
rect 499 593 533 595
rect 499 521 533 527
rect 499 449 533 459
rect 499 377 533 391
rect 499 305 533 323
rect 499 233 533 255
rect 499 161 533 187
rect 499 89 533 119
rect 499 17 533 51
rect 499 -51 533 -17
rect 499 -119 533 -89
rect 499 -187 533 -161
rect 499 -255 533 -233
rect 499 -323 533 -305
rect 499 -391 533 -377
rect 499 -459 533 -449
rect 499 -527 533 -521
rect 499 -595 533 -593
rect 499 -631 533 -629
rect 499 -703 533 -697
rect 499 -775 533 -765
rect 499 -847 533 -833
rect 499 -919 533 -901
rect 499 -991 533 -969
rect 499 -1063 533 -1037
rect 499 -1135 533 -1105
rect 499 -1207 533 -1173
rect 499 -1275 533 -1241
rect 499 -1343 533 -1313
rect 499 -1411 533 -1385
rect 499 -1479 533 -1457
rect 499 -1547 533 -1529
rect 499 -1615 533 -1601
rect 499 -1683 533 -1673
rect 499 -1751 533 -1745
rect 499 -1819 533 -1817
rect 499 -1855 533 -1853
rect 499 -1927 533 -1921
rect 499 -1999 533 -1989
rect 499 -2071 533 -2057
rect 499 -2143 533 -2125
rect 499 -2215 533 -2193
rect 499 -2287 533 -2261
rect 499 -2359 533 -2329
rect 499 -2431 533 -2397
rect 499 -2504 533 -2465
rect 757 2465 791 2504
rect 757 2397 791 2431
rect 757 2329 791 2359
rect 757 2261 791 2287
rect 757 2193 791 2215
rect 757 2125 791 2143
rect 757 2057 791 2071
rect 757 1989 791 1999
rect 757 1921 791 1927
rect 757 1853 791 1855
rect 757 1817 791 1819
rect 757 1745 791 1751
rect 757 1673 791 1683
rect 757 1601 791 1615
rect 757 1529 791 1547
rect 757 1457 791 1479
rect 757 1385 791 1411
rect 757 1313 791 1343
rect 757 1241 791 1275
rect 757 1173 791 1207
rect 757 1105 791 1135
rect 757 1037 791 1063
rect 757 969 791 991
rect 757 901 791 919
rect 757 833 791 847
rect 757 765 791 775
rect 757 697 791 703
rect 757 629 791 631
rect 757 593 791 595
rect 757 521 791 527
rect 757 449 791 459
rect 757 377 791 391
rect 757 305 791 323
rect 757 233 791 255
rect 757 161 791 187
rect 757 89 791 119
rect 757 17 791 51
rect 757 -51 791 -17
rect 757 -119 791 -89
rect 757 -187 791 -161
rect 757 -255 791 -233
rect 757 -323 791 -305
rect 757 -391 791 -377
rect 757 -459 791 -449
rect 757 -527 791 -521
rect 757 -595 791 -593
rect 757 -631 791 -629
rect 757 -703 791 -697
rect 757 -775 791 -765
rect 757 -847 791 -833
rect 757 -919 791 -901
rect 757 -991 791 -969
rect 757 -1063 791 -1037
rect 757 -1135 791 -1105
rect 757 -1207 791 -1173
rect 757 -1275 791 -1241
rect 757 -1343 791 -1313
rect 757 -1411 791 -1385
rect 757 -1479 791 -1457
rect 757 -1547 791 -1529
rect 757 -1615 791 -1601
rect 757 -1683 791 -1673
rect 757 -1751 791 -1745
rect 757 -1819 791 -1817
rect 757 -1855 791 -1853
rect 757 -1927 791 -1921
rect 757 -1999 791 -1989
rect 757 -2071 791 -2057
rect 757 -2143 791 -2125
rect 757 -2215 791 -2193
rect 757 -2287 791 -2261
rect 757 -2359 791 -2329
rect 757 -2431 791 -2397
rect 757 -2504 791 -2465
rect 1015 2465 1049 2504
rect 1015 2397 1049 2431
rect 1015 2329 1049 2359
rect 1015 2261 1049 2287
rect 1015 2193 1049 2215
rect 1015 2125 1049 2143
rect 1015 2057 1049 2071
rect 1015 1989 1049 1999
rect 1015 1921 1049 1927
rect 1015 1853 1049 1855
rect 1015 1817 1049 1819
rect 1015 1745 1049 1751
rect 1015 1673 1049 1683
rect 1015 1601 1049 1615
rect 1015 1529 1049 1547
rect 1015 1457 1049 1479
rect 1015 1385 1049 1411
rect 1015 1313 1049 1343
rect 1015 1241 1049 1275
rect 1015 1173 1049 1207
rect 1015 1105 1049 1135
rect 1015 1037 1049 1063
rect 1015 969 1049 991
rect 1015 901 1049 919
rect 1015 833 1049 847
rect 1015 765 1049 775
rect 1015 697 1049 703
rect 1015 629 1049 631
rect 1015 593 1049 595
rect 1015 521 1049 527
rect 1015 449 1049 459
rect 1015 377 1049 391
rect 1015 305 1049 323
rect 1015 233 1049 255
rect 1015 161 1049 187
rect 1015 89 1049 119
rect 1015 17 1049 51
rect 1015 -51 1049 -17
rect 1015 -119 1049 -89
rect 1015 -187 1049 -161
rect 1015 -255 1049 -233
rect 1015 -323 1049 -305
rect 1015 -391 1049 -377
rect 1015 -459 1049 -449
rect 1015 -527 1049 -521
rect 1015 -595 1049 -593
rect 1015 -631 1049 -629
rect 1015 -703 1049 -697
rect 1015 -775 1049 -765
rect 1015 -847 1049 -833
rect 1015 -919 1049 -901
rect 1015 -991 1049 -969
rect 1015 -1063 1049 -1037
rect 1015 -1135 1049 -1105
rect 1015 -1207 1049 -1173
rect 1015 -1275 1049 -1241
rect 1015 -1343 1049 -1313
rect 1015 -1411 1049 -1385
rect 1015 -1479 1049 -1457
rect 1015 -1547 1049 -1529
rect 1015 -1615 1049 -1601
rect 1015 -1683 1049 -1673
rect 1015 -1751 1049 -1745
rect 1015 -1819 1049 -1817
rect 1015 -1855 1049 -1853
rect 1015 -1927 1049 -1921
rect 1015 -1999 1049 -1989
rect 1015 -2071 1049 -2057
rect 1015 -2143 1049 -2125
rect 1015 -2215 1049 -2193
rect 1015 -2287 1049 -2261
rect 1015 -2359 1049 -2329
rect 1015 -2431 1049 -2397
rect 1015 -2504 1049 -2465
rect 1273 2465 1307 2504
rect 1273 2397 1307 2431
rect 1273 2329 1307 2359
rect 1273 2261 1307 2287
rect 1273 2193 1307 2215
rect 1273 2125 1307 2143
rect 1273 2057 1307 2071
rect 1273 1989 1307 1999
rect 1273 1921 1307 1927
rect 1273 1853 1307 1855
rect 1273 1817 1307 1819
rect 1273 1745 1307 1751
rect 1273 1673 1307 1683
rect 1273 1601 1307 1615
rect 1273 1529 1307 1547
rect 1273 1457 1307 1479
rect 1273 1385 1307 1411
rect 1273 1313 1307 1343
rect 1273 1241 1307 1275
rect 1273 1173 1307 1207
rect 1273 1105 1307 1135
rect 1273 1037 1307 1063
rect 1273 969 1307 991
rect 1273 901 1307 919
rect 1273 833 1307 847
rect 1273 765 1307 775
rect 1273 697 1307 703
rect 1273 629 1307 631
rect 1273 593 1307 595
rect 1273 521 1307 527
rect 1273 449 1307 459
rect 1273 377 1307 391
rect 1273 305 1307 323
rect 1273 233 1307 255
rect 1273 161 1307 187
rect 1273 89 1307 119
rect 1273 17 1307 51
rect 1273 -51 1307 -17
rect 1273 -119 1307 -89
rect 1273 -187 1307 -161
rect 1273 -255 1307 -233
rect 1273 -323 1307 -305
rect 1273 -391 1307 -377
rect 1273 -459 1307 -449
rect 1273 -527 1307 -521
rect 1273 -595 1307 -593
rect 1273 -631 1307 -629
rect 1273 -703 1307 -697
rect 1273 -775 1307 -765
rect 1273 -847 1307 -833
rect 1273 -919 1307 -901
rect 1273 -991 1307 -969
rect 1273 -1063 1307 -1037
rect 1273 -1135 1307 -1105
rect 1273 -1207 1307 -1173
rect 1273 -1275 1307 -1241
rect 1273 -1343 1307 -1313
rect 1273 -1411 1307 -1385
rect 1273 -1479 1307 -1457
rect 1273 -1547 1307 -1529
rect 1273 -1615 1307 -1601
rect 1273 -1683 1307 -1673
rect 1273 -1751 1307 -1745
rect 1273 -1819 1307 -1817
rect 1273 -1855 1307 -1853
rect 1273 -1927 1307 -1921
rect 1273 -1999 1307 -1989
rect 1273 -2071 1307 -2057
rect 1273 -2143 1307 -2125
rect 1273 -2215 1307 -2193
rect 1273 -2287 1307 -2261
rect 1273 -2359 1307 -2329
rect 1273 -2431 1307 -2397
rect 1273 -2504 1307 -2465
rect 1387 2499 1421 2533
rect 1387 2431 1421 2465
rect 1387 2363 1421 2397
rect 1387 2295 1421 2329
rect 1387 2227 1421 2261
rect 1387 2159 1421 2193
rect 1387 2091 1421 2125
rect 1387 2023 1421 2057
rect 1387 1955 1421 1989
rect 1387 1887 1421 1921
rect 1387 1819 1421 1853
rect 1387 1751 1421 1785
rect 1387 1683 1421 1717
rect 1387 1615 1421 1649
rect 1387 1547 1421 1581
rect 1387 1479 1421 1513
rect 1387 1411 1421 1445
rect 1387 1343 1421 1377
rect 1387 1275 1421 1309
rect 1387 1207 1421 1241
rect 1387 1139 1421 1173
rect 1387 1071 1421 1105
rect 1387 1003 1421 1037
rect 1387 935 1421 969
rect 1387 867 1421 901
rect 1387 799 1421 833
rect 1387 731 1421 765
rect 1387 663 1421 697
rect 1387 595 1421 629
rect 1387 527 1421 561
rect 1387 459 1421 493
rect 1387 391 1421 425
rect 1387 323 1421 357
rect 1387 255 1421 289
rect 1387 187 1421 221
rect 1387 119 1421 153
rect 1387 51 1421 85
rect 1387 -17 1421 17
rect 1387 -85 1421 -51
rect 1387 -153 1421 -119
rect 1387 -221 1421 -187
rect 1387 -289 1421 -255
rect 1387 -357 1421 -323
rect 1387 -425 1421 -391
rect 1387 -493 1421 -459
rect 1387 -561 1421 -527
rect 1387 -629 1421 -595
rect 1387 -697 1421 -663
rect 1387 -765 1421 -731
rect 1387 -833 1421 -799
rect 1387 -901 1421 -867
rect 1387 -969 1421 -935
rect 1387 -1037 1421 -1003
rect 1387 -1105 1421 -1071
rect 1387 -1173 1421 -1139
rect 1387 -1241 1421 -1207
rect 1387 -1309 1421 -1275
rect 1387 -1377 1421 -1343
rect 1387 -1445 1421 -1411
rect 1387 -1513 1421 -1479
rect 1387 -1581 1421 -1547
rect 1387 -1649 1421 -1615
rect 1387 -1717 1421 -1683
rect 1387 -1785 1421 -1751
rect 1387 -1853 1421 -1819
rect 1387 -1921 1421 -1887
rect 1387 -1989 1421 -1955
rect 1387 -2057 1421 -2023
rect 1387 -2125 1421 -2091
rect 1387 -2193 1421 -2159
rect 1387 -2261 1421 -2227
rect 1387 -2329 1421 -2295
rect 1387 -2397 1421 -2363
rect 1387 -2465 1421 -2431
rect 1387 -2533 1421 -2499
rect -1421 -2640 -1387 -2567
rect -1261 -2572 -1214 -2538
rect -1178 -2572 -1144 -2538
rect -1108 -2572 -1061 -2538
rect -1003 -2572 -956 -2538
rect -920 -2572 -886 -2538
rect -850 -2572 -803 -2538
rect -745 -2572 -698 -2538
rect -662 -2572 -628 -2538
rect -592 -2572 -545 -2538
rect -487 -2572 -440 -2538
rect -404 -2572 -370 -2538
rect -334 -2572 -287 -2538
rect -229 -2572 -182 -2538
rect -146 -2572 -112 -2538
rect -76 -2572 -29 -2538
rect 29 -2572 76 -2538
rect 112 -2572 146 -2538
rect 182 -2572 229 -2538
rect 287 -2572 334 -2538
rect 370 -2572 404 -2538
rect 440 -2572 487 -2538
rect 545 -2572 592 -2538
rect 628 -2572 662 -2538
rect 698 -2572 745 -2538
rect 803 -2572 850 -2538
rect 886 -2572 920 -2538
rect 956 -2572 1003 -2538
rect 1061 -2572 1108 -2538
rect 1144 -2572 1178 -2538
rect 1214 -2572 1261 -2538
rect 1387 -2640 1421 -2567
rect -1421 -2674 -1309 -2640
rect -1275 -2674 -1241 -2640
rect -1207 -2674 -1173 -2640
rect -1139 -2674 -1105 -2640
rect -1071 -2674 -1037 -2640
rect -1003 -2674 -969 -2640
rect -935 -2674 -901 -2640
rect -867 -2674 -833 -2640
rect -799 -2674 -765 -2640
rect -731 -2674 -697 -2640
rect -663 -2674 -629 -2640
rect -595 -2674 -561 -2640
rect -527 -2674 -493 -2640
rect -459 -2674 -425 -2640
rect -391 -2674 -357 -2640
rect -323 -2674 -289 -2640
rect -255 -2674 -221 -2640
rect -187 -2674 -153 -2640
rect -119 -2674 -85 -2640
rect -51 -2674 -17 -2640
rect 17 -2674 51 -2640
rect 85 -2674 119 -2640
rect 153 -2674 187 -2640
rect 221 -2674 255 -2640
rect 289 -2674 323 -2640
rect 357 -2674 391 -2640
rect 425 -2674 459 -2640
rect 493 -2674 527 -2640
rect 561 -2674 595 -2640
rect 629 -2674 663 -2640
rect 697 -2674 731 -2640
rect 765 -2674 799 -2640
rect 833 -2674 867 -2640
rect 901 -2674 935 -2640
rect 969 -2674 1003 -2640
rect 1037 -2674 1071 -2640
rect 1105 -2674 1139 -2640
rect 1173 -2674 1207 -2640
rect 1241 -2674 1275 -2640
rect 1309 -2674 1421 -2640
<< viali >>
rect -1214 2538 -1212 2572
rect -1212 2538 -1180 2572
rect -1142 2538 -1110 2572
rect -1110 2538 -1108 2572
rect -956 2538 -954 2572
rect -954 2538 -922 2572
rect -884 2538 -852 2572
rect -852 2538 -850 2572
rect -698 2538 -696 2572
rect -696 2538 -664 2572
rect -626 2538 -594 2572
rect -594 2538 -592 2572
rect -440 2538 -438 2572
rect -438 2538 -406 2572
rect -368 2538 -336 2572
rect -336 2538 -334 2572
rect -182 2538 -180 2572
rect -180 2538 -148 2572
rect -110 2538 -78 2572
rect -78 2538 -76 2572
rect 76 2538 78 2572
rect 78 2538 110 2572
rect 148 2538 180 2572
rect 180 2538 182 2572
rect 334 2538 336 2572
rect 336 2538 368 2572
rect 406 2538 438 2572
rect 438 2538 440 2572
rect 592 2538 594 2572
rect 594 2538 626 2572
rect 664 2538 696 2572
rect 696 2538 698 2572
rect 850 2538 852 2572
rect 852 2538 884 2572
rect 922 2538 954 2572
rect 954 2538 956 2572
rect 1108 2538 1110 2572
rect 1110 2538 1142 2572
rect 1180 2538 1212 2572
rect 1212 2538 1214 2572
rect -1307 2431 -1273 2465
rect -1307 2363 -1273 2393
rect -1307 2359 -1273 2363
rect -1307 2295 -1273 2321
rect -1307 2287 -1273 2295
rect -1307 2227 -1273 2249
rect -1307 2215 -1273 2227
rect -1307 2159 -1273 2177
rect -1307 2143 -1273 2159
rect -1307 2091 -1273 2105
rect -1307 2071 -1273 2091
rect -1307 2023 -1273 2033
rect -1307 1999 -1273 2023
rect -1307 1955 -1273 1961
rect -1307 1927 -1273 1955
rect -1307 1887 -1273 1889
rect -1307 1855 -1273 1887
rect -1307 1785 -1273 1817
rect -1307 1783 -1273 1785
rect -1307 1717 -1273 1745
rect -1307 1711 -1273 1717
rect -1307 1649 -1273 1673
rect -1307 1639 -1273 1649
rect -1307 1581 -1273 1601
rect -1307 1567 -1273 1581
rect -1307 1513 -1273 1529
rect -1307 1495 -1273 1513
rect -1307 1445 -1273 1457
rect -1307 1423 -1273 1445
rect -1307 1377 -1273 1385
rect -1307 1351 -1273 1377
rect -1307 1309 -1273 1313
rect -1307 1279 -1273 1309
rect -1307 1207 -1273 1241
rect -1307 1139 -1273 1169
rect -1307 1135 -1273 1139
rect -1307 1071 -1273 1097
rect -1307 1063 -1273 1071
rect -1307 1003 -1273 1025
rect -1307 991 -1273 1003
rect -1307 935 -1273 953
rect -1307 919 -1273 935
rect -1307 867 -1273 881
rect -1307 847 -1273 867
rect -1307 799 -1273 809
rect -1307 775 -1273 799
rect -1307 731 -1273 737
rect -1307 703 -1273 731
rect -1307 663 -1273 665
rect -1307 631 -1273 663
rect -1307 561 -1273 593
rect -1307 559 -1273 561
rect -1307 493 -1273 521
rect -1307 487 -1273 493
rect -1307 425 -1273 449
rect -1307 415 -1273 425
rect -1307 357 -1273 377
rect -1307 343 -1273 357
rect -1307 289 -1273 305
rect -1307 271 -1273 289
rect -1307 221 -1273 233
rect -1307 199 -1273 221
rect -1307 153 -1273 161
rect -1307 127 -1273 153
rect -1307 85 -1273 89
rect -1307 55 -1273 85
rect -1307 -17 -1273 17
rect -1307 -85 -1273 -55
rect -1307 -89 -1273 -85
rect -1307 -153 -1273 -127
rect -1307 -161 -1273 -153
rect -1307 -221 -1273 -199
rect -1307 -233 -1273 -221
rect -1307 -289 -1273 -271
rect -1307 -305 -1273 -289
rect -1307 -357 -1273 -343
rect -1307 -377 -1273 -357
rect -1307 -425 -1273 -415
rect -1307 -449 -1273 -425
rect -1307 -493 -1273 -487
rect -1307 -521 -1273 -493
rect -1307 -561 -1273 -559
rect -1307 -593 -1273 -561
rect -1307 -663 -1273 -631
rect -1307 -665 -1273 -663
rect -1307 -731 -1273 -703
rect -1307 -737 -1273 -731
rect -1307 -799 -1273 -775
rect -1307 -809 -1273 -799
rect -1307 -867 -1273 -847
rect -1307 -881 -1273 -867
rect -1307 -935 -1273 -919
rect -1307 -953 -1273 -935
rect -1307 -1003 -1273 -991
rect -1307 -1025 -1273 -1003
rect -1307 -1071 -1273 -1063
rect -1307 -1097 -1273 -1071
rect -1307 -1139 -1273 -1135
rect -1307 -1169 -1273 -1139
rect -1307 -1241 -1273 -1207
rect -1307 -1309 -1273 -1279
rect -1307 -1313 -1273 -1309
rect -1307 -1377 -1273 -1351
rect -1307 -1385 -1273 -1377
rect -1307 -1445 -1273 -1423
rect -1307 -1457 -1273 -1445
rect -1307 -1513 -1273 -1495
rect -1307 -1529 -1273 -1513
rect -1307 -1581 -1273 -1567
rect -1307 -1601 -1273 -1581
rect -1307 -1649 -1273 -1639
rect -1307 -1673 -1273 -1649
rect -1307 -1717 -1273 -1711
rect -1307 -1745 -1273 -1717
rect -1307 -1785 -1273 -1783
rect -1307 -1817 -1273 -1785
rect -1307 -1887 -1273 -1855
rect -1307 -1889 -1273 -1887
rect -1307 -1955 -1273 -1927
rect -1307 -1961 -1273 -1955
rect -1307 -2023 -1273 -1999
rect -1307 -2033 -1273 -2023
rect -1307 -2091 -1273 -2071
rect -1307 -2105 -1273 -2091
rect -1307 -2159 -1273 -2143
rect -1307 -2177 -1273 -2159
rect -1307 -2227 -1273 -2215
rect -1307 -2249 -1273 -2227
rect -1307 -2295 -1273 -2287
rect -1307 -2321 -1273 -2295
rect -1307 -2363 -1273 -2359
rect -1307 -2393 -1273 -2363
rect -1307 -2465 -1273 -2431
rect -1049 2431 -1015 2465
rect -1049 2363 -1015 2393
rect -1049 2359 -1015 2363
rect -1049 2295 -1015 2321
rect -1049 2287 -1015 2295
rect -1049 2227 -1015 2249
rect -1049 2215 -1015 2227
rect -1049 2159 -1015 2177
rect -1049 2143 -1015 2159
rect -1049 2091 -1015 2105
rect -1049 2071 -1015 2091
rect -1049 2023 -1015 2033
rect -1049 1999 -1015 2023
rect -1049 1955 -1015 1961
rect -1049 1927 -1015 1955
rect -1049 1887 -1015 1889
rect -1049 1855 -1015 1887
rect -1049 1785 -1015 1817
rect -1049 1783 -1015 1785
rect -1049 1717 -1015 1745
rect -1049 1711 -1015 1717
rect -1049 1649 -1015 1673
rect -1049 1639 -1015 1649
rect -1049 1581 -1015 1601
rect -1049 1567 -1015 1581
rect -1049 1513 -1015 1529
rect -1049 1495 -1015 1513
rect -1049 1445 -1015 1457
rect -1049 1423 -1015 1445
rect -1049 1377 -1015 1385
rect -1049 1351 -1015 1377
rect -1049 1309 -1015 1313
rect -1049 1279 -1015 1309
rect -1049 1207 -1015 1241
rect -1049 1139 -1015 1169
rect -1049 1135 -1015 1139
rect -1049 1071 -1015 1097
rect -1049 1063 -1015 1071
rect -1049 1003 -1015 1025
rect -1049 991 -1015 1003
rect -1049 935 -1015 953
rect -1049 919 -1015 935
rect -1049 867 -1015 881
rect -1049 847 -1015 867
rect -1049 799 -1015 809
rect -1049 775 -1015 799
rect -1049 731 -1015 737
rect -1049 703 -1015 731
rect -1049 663 -1015 665
rect -1049 631 -1015 663
rect -1049 561 -1015 593
rect -1049 559 -1015 561
rect -1049 493 -1015 521
rect -1049 487 -1015 493
rect -1049 425 -1015 449
rect -1049 415 -1015 425
rect -1049 357 -1015 377
rect -1049 343 -1015 357
rect -1049 289 -1015 305
rect -1049 271 -1015 289
rect -1049 221 -1015 233
rect -1049 199 -1015 221
rect -1049 153 -1015 161
rect -1049 127 -1015 153
rect -1049 85 -1015 89
rect -1049 55 -1015 85
rect -1049 -17 -1015 17
rect -1049 -85 -1015 -55
rect -1049 -89 -1015 -85
rect -1049 -153 -1015 -127
rect -1049 -161 -1015 -153
rect -1049 -221 -1015 -199
rect -1049 -233 -1015 -221
rect -1049 -289 -1015 -271
rect -1049 -305 -1015 -289
rect -1049 -357 -1015 -343
rect -1049 -377 -1015 -357
rect -1049 -425 -1015 -415
rect -1049 -449 -1015 -425
rect -1049 -493 -1015 -487
rect -1049 -521 -1015 -493
rect -1049 -561 -1015 -559
rect -1049 -593 -1015 -561
rect -1049 -663 -1015 -631
rect -1049 -665 -1015 -663
rect -1049 -731 -1015 -703
rect -1049 -737 -1015 -731
rect -1049 -799 -1015 -775
rect -1049 -809 -1015 -799
rect -1049 -867 -1015 -847
rect -1049 -881 -1015 -867
rect -1049 -935 -1015 -919
rect -1049 -953 -1015 -935
rect -1049 -1003 -1015 -991
rect -1049 -1025 -1015 -1003
rect -1049 -1071 -1015 -1063
rect -1049 -1097 -1015 -1071
rect -1049 -1139 -1015 -1135
rect -1049 -1169 -1015 -1139
rect -1049 -1241 -1015 -1207
rect -1049 -1309 -1015 -1279
rect -1049 -1313 -1015 -1309
rect -1049 -1377 -1015 -1351
rect -1049 -1385 -1015 -1377
rect -1049 -1445 -1015 -1423
rect -1049 -1457 -1015 -1445
rect -1049 -1513 -1015 -1495
rect -1049 -1529 -1015 -1513
rect -1049 -1581 -1015 -1567
rect -1049 -1601 -1015 -1581
rect -1049 -1649 -1015 -1639
rect -1049 -1673 -1015 -1649
rect -1049 -1717 -1015 -1711
rect -1049 -1745 -1015 -1717
rect -1049 -1785 -1015 -1783
rect -1049 -1817 -1015 -1785
rect -1049 -1887 -1015 -1855
rect -1049 -1889 -1015 -1887
rect -1049 -1955 -1015 -1927
rect -1049 -1961 -1015 -1955
rect -1049 -2023 -1015 -1999
rect -1049 -2033 -1015 -2023
rect -1049 -2091 -1015 -2071
rect -1049 -2105 -1015 -2091
rect -1049 -2159 -1015 -2143
rect -1049 -2177 -1015 -2159
rect -1049 -2227 -1015 -2215
rect -1049 -2249 -1015 -2227
rect -1049 -2295 -1015 -2287
rect -1049 -2321 -1015 -2295
rect -1049 -2363 -1015 -2359
rect -1049 -2393 -1015 -2363
rect -1049 -2465 -1015 -2431
rect -791 2431 -757 2465
rect -791 2363 -757 2393
rect -791 2359 -757 2363
rect -791 2295 -757 2321
rect -791 2287 -757 2295
rect -791 2227 -757 2249
rect -791 2215 -757 2227
rect -791 2159 -757 2177
rect -791 2143 -757 2159
rect -791 2091 -757 2105
rect -791 2071 -757 2091
rect -791 2023 -757 2033
rect -791 1999 -757 2023
rect -791 1955 -757 1961
rect -791 1927 -757 1955
rect -791 1887 -757 1889
rect -791 1855 -757 1887
rect -791 1785 -757 1817
rect -791 1783 -757 1785
rect -791 1717 -757 1745
rect -791 1711 -757 1717
rect -791 1649 -757 1673
rect -791 1639 -757 1649
rect -791 1581 -757 1601
rect -791 1567 -757 1581
rect -791 1513 -757 1529
rect -791 1495 -757 1513
rect -791 1445 -757 1457
rect -791 1423 -757 1445
rect -791 1377 -757 1385
rect -791 1351 -757 1377
rect -791 1309 -757 1313
rect -791 1279 -757 1309
rect -791 1207 -757 1241
rect -791 1139 -757 1169
rect -791 1135 -757 1139
rect -791 1071 -757 1097
rect -791 1063 -757 1071
rect -791 1003 -757 1025
rect -791 991 -757 1003
rect -791 935 -757 953
rect -791 919 -757 935
rect -791 867 -757 881
rect -791 847 -757 867
rect -791 799 -757 809
rect -791 775 -757 799
rect -791 731 -757 737
rect -791 703 -757 731
rect -791 663 -757 665
rect -791 631 -757 663
rect -791 561 -757 593
rect -791 559 -757 561
rect -791 493 -757 521
rect -791 487 -757 493
rect -791 425 -757 449
rect -791 415 -757 425
rect -791 357 -757 377
rect -791 343 -757 357
rect -791 289 -757 305
rect -791 271 -757 289
rect -791 221 -757 233
rect -791 199 -757 221
rect -791 153 -757 161
rect -791 127 -757 153
rect -791 85 -757 89
rect -791 55 -757 85
rect -791 -17 -757 17
rect -791 -85 -757 -55
rect -791 -89 -757 -85
rect -791 -153 -757 -127
rect -791 -161 -757 -153
rect -791 -221 -757 -199
rect -791 -233 -757 -221
rect -791 -289 -757 -271
rect -791 -305 -757 -289
rect -791 -357 -757 -343
rect -791 -377 -757 -357
rect -791 -425 -757 -415
rect -791 -449 -757 -425
rect -791 -493 -757 -487
rect -791 -521 -757 -493
rect -791 -561 -757 -559
rect -791 -593 -757 -561
rect -791 -663 -757 -631
rect -791 -665 -757 -663
rect -791 -731 -757 -703
rect -791 -737 -757 -731
rect -791 -799 -757 -775
rect -791 -809 -757 -799
rect -791 -867 -757 -847
rect -791 -881 -757 -867
rect -791 -935 -757 -919
rect -791 -953 -757 -935
rect -791 -1003 -757 -991
rect -791 -1025 -757 -1003
rect -791 -1071 -757 -1063
rect -791 -1097 -757 -1071
rect -791 -1139 -757 -1135
rect -791 -1169 -757 -1139
rect -791 -1241 -757 -1207
rect -791 -1309 -757 -1279
rect -791 -1313 -757 -1309
rect -791 -1377 -757 -1351
rect -791 -1385 -757 -1377
rect -791 -1445 -757 -1423
rect -791 -1457 -757 -1445
rect -791 -1513 -757 -1495
rect -791 -1529 -757 -1513
rect -791 -1581 -757 -1567
rect -791 -1601 -757 -1581
rect -791 -1649 -757 -1639
rect -791 -1673 -757 -1649
rect -791 -1717 -757 -1711
rect -791 -1745 -757 -1717
rect -791 -1785 -757 -1783
rect -791 -1817 -757 -1785
rect -791 -1887 -757 -1855
rect -791 -1889 -757 -1887
rect -791 -1955 -757 -1927
rect -791 -1961 -757 -1955
rect -791 -2023 -757 -1999
rect -791 -2033 -757 -2023
rect -791 -2091 -757 -2071
rect -791 -2105 -757 -2091
rect -791 -2159 -757 -2143
rect -791 -2177 -757 -2159
rect -791 -2227 -757 -2215
rect -791 -2249 -757 -2227
rect -791 -2295 -757 -2287
rect -791 -2321 -757 -2295
rect -791 -2363 -757 -2359
rect -791 -2393 -757 -2363
rect -791 -2465 -757 -2431
rect -533 2431 -499 2465
rect -533 2363 -499 2393
rect -533 2359 -499 2363
rect -533 2295 -499 2321
rect -533 2287 -499 2295
rect -533 2227 -499 2249
rect -533 2215 -499 2227
rect -533 2159 -499 2177
rect -533 2143 -499 2159
rect -533 2091 -499 2105
rect -533 2071 -499 2091
rect -533 2023 -499 2033
rect -533 1999 -499 2023
rect -533 1955 -499 1961
rect -533 1927 -499 1955
rect -533 1887 -499 1889
rect -533 1855 -499 1887
rect -533 1785 -499 1817
rect -533 1783 -499 1785
rect -533 1717 -499 1745
rect -533 1711 -499 1717
rect -533 1649 -499 1673
rect -533 1639 -499 1649
rect -533 1581 -499 1601
rect -533 1567 -499 1581
rect -533 1513 -499 1529
rect -533 1495 -499 1513
rect -533 1445 -499 1457
rect -533 1423 -499 1445
rect -533 1377 -499 1385
rect -533 1351 -499 1377
rect -533 1309 -499 1313
rect -533 1279 -499 1309
rect -533 1207 -499 1241
rect -533 1139 -499 1169
rect -533 1135 -499 1139
rect -533 1071 -499 1097
rect -533 1063 -499 1071
rect -533 1003 -499 1025
rect -533 991 -499 1003
rect -533 935 -499 953
rect -533 919 -499 935
rect -533 867 -499 881
rect -533 847 -499 867
rect -533 799 -499 809
rect -533 775 -499 799
rect -533 731 -499 737
rect -533 703 -499 731
rect -533 663 -499 665
rect -533 631 -499 663
rect -533 561 -499 593
rect -533 559 -499 561
rect -533 493 -499 521
rect -533 487 -499 493
rect -533 425 -499 449
rect -533 415 -499 425
rect -533 357 -499 377
rect -533 343 -499 357
rect -533 289 -499 305
rect -533 271 -499 289
rect -533 221 -499 233
rect -533 199 -499 221
rect -533 153 -499 161
rect -533 127 -499 153
rect -533 85 -499 89
rect -533 55 -499 85
rect -533 -17 -499 17
rect -533 -85 -499 -55
rect -533 -89 -499 -85
rect -533 -153 -499 -127
rect -533 -161 -499 -153
rect -533 -221 -499 -199
rect -533 -233 -499 -221
rect -533 -289 -499 -271
rect -533 -305 -499 -289
rect -533 -357 -499 -343
rect -533 -377 -499 -357
rect -533 -425 -499 -415
rect -533 -449 -499 -425
rect -533 -493 -499 -487
rect -533 -521 -499 -493
rect -533 -561 -499 -559
rect -533 -593 -499 -561
rect -533 -663 -499 -631
rect -533 -665 -499 -663
rect -533 -731 -499 -703
rect -533 -737 -499 -731
rect -533 -799 -499 -775
rect -533 -809 -499 -799
rect -533 -867 -499 -847
rect -533 -881 -499 -867
rect -533 -935 -499 -919
rect -533 -953 -499 -935
rect -533 -1003 -499 -991
rect -533 -1025 -499 -1003
rect -533 -1071 -499 -1063
rect -533 -1097 -499 -1071
rect -533 -1139 -499 -1135
rect -533 -1169 -499 -1139
rect -533 -1241 -499 -1207
rect -533 -1309 -499 -1279
rect -533 -1313 -499 -1309
rect -533 -1377 -499 -1351
rect -533 -1385 -499 -1377
rect -533 -1445 -499 -1423
rect -533 -1457 -499 -1445
rect -533 -1513 -499 -1495
rect -533 -1529 -499 -1513
rect -533 -1581 -499 -1567
rect -533 -1601 -499 -1581
rect -533 -1649 -499 -1639
rect -533 -1673 -499 -1649
rect -533 -1717 -499 -1711
rect -533 -1745 -499 -1717
rect -533 -1785 -499 -1783
rect -533 -1817 -499 -1785
rect -533 -1887 -499 -1855
rect -533 -1889 -499 -1887
rect -533 -1955 -499 -1927
rect -533 -1961 -499 -1955
rect -533 -2023 -499 -1999
rect -533 -2033 -499 -2023
rect -533 -2091 -499 -2071
rect -533 -2105 -499 -2091
rect -533 -2159 -499 -2143
rect -533 -2177 -499 -2159
rect -533 -2227 -499 -2215
rect -533 -2249 -499 -2227
rect -533 -2295 -499 -2287
rect -533 -2321 -499 -2295
rect -533 -2363 -499 -2359
rect -533 -2393 -499 -2363
rect -533 -2465 -499 -2431
rect -275 2431 -241 2465
rect -275 2363 -241 2393
rect -275 2359 -241 2363
rect -275 2295 -241 2321
rect -275 2287 -241 2295
rect -275 2227 -241 2249
rect -275 2215 -241 2227
rect -275 2159 -241 2177
rect -275 2143 -241 2159
rect -275 2091 -241 2105
rect -275 2071 -241 2091
rect -275 2023 -241 2033
rect -275 1999 -241 2023
rect -275 1955 -241 1961
rect -275 1927 -241 1955
rect -275 1887 -241 1889
rect -275 1855 -241 1887
rect -275 1785 -241 1817
rect -275 1783 -241 1785
rect -275 1717 -241 1745
rect -275 1711 -241 1717
rect -275 1649 -241 1673
rect -275 1639 -241 1649
rect -275 1581 -241 1601
rect -275 1567 -241 1581
rect -275 1513 -241 1529
rect -275 1495 -241 1513
rect -275 1445 -241 1457
rect -275 1423 -241 1445
rect -275 1377 -241 1385
rect -275 1351 -241 1377
rect -275 1309 -241 1313
rect -275 1279 -241 1309
rect -275 1207 -241 1241
rect -275 1139 -241 1169
rect -275 1135 -241 1139
rect -275 1071 -241 1097
rect -275 1063 -241 1071
rect -275 1003 -241 1025
rect -275 991 -241 1003
rect -275 935 -241 953
rect -275 919 -241 935
rect -275 867 -241 881
rect -275 847 -241 867
rect -275 799 -241 809
rect -275 775 -241 799
rect -275 731 -241 737
rect -275 703 -241 731
rect -275 663 -241 665
rect -275 631 -241 663
rect -275 561 -241 593
rect -275 559 -241 561
rect -275 493 -241 521
rect -275 487 -241 493
rect -275 425 -241 449
rect -275 415 -241 425
rect -275 357 -241 377
rect -275 343 -241 357
rect -275 289 -241 305
rect -275 271 -241 289
rect -275 221 -241 233
rect -275 199 -241 221
rect -275 153 -241 161
rect -275 127 -241 153
rect -275 85 -241 89
rect -275 55 -241 85
rect -275 -17 -241 17
rect -275 -85 -241 -55
rect -275 -89 -241 -85
rect -275 -153 -241 -127
rect -275 -161 -241 -153
rect -275 -221 -241 -199
rect -275 -233 -241 -221
rect -275 -289 -241 -271
rect -275 -305 -241 -289
rect -275 -357 -241 -343
rect -275 -377 -241 -357
rect -275 -425 -241 -415
rect -275 -449 -241 -425
rect -275 -493 -241 -487
rect -275 -521 -241 -493
rect -275 -561 -241 -559
rect -275 -593 -241 -561
rect -275 -663 -241 -631
rect -275 -665 -241 -663
rect -275 -731 -241 -703
rect -275 -737 -241 -731
rect -275 -799 -241 -775
rect -275 -809 -241 -799
rect -275 -867 -241 -847
rect -275 -881 -241 -867
rect -275 -935 -241 -919
rect -275 -953 -241 -935
rect -275 -1003 -241 -991
rect -275 -1025 -241 -1003
rect -275 -1071 -241 -1063
rect -275 -1097 -241 -1071
rect -275 -1139 -241 -1135
rect -275 -1169 -241 -1139
rect -275 -1241 -241 -1207
rect -275 -1309 -241 -1279
rect -275 -1313 -241 -1309
rect -275 -1377 -241 -1351
rect -275 -1385 -241 -1377
rect -275 -1445 -241 -1423
rect -275 -1457 -241 -1445
rect -275 -1513 -241 -1495
rect -275 -1529 -241 -1513
rect -275 -1581 -241 -1567
rect -275 -1601 -241 -1581
rect -275 -1649 -241 -1639
rect -275 -1673 -241 -1649
rect -275 -1717 -241 -1711
rect -275 -1745 -241 -1717
rect -275 -1785 -241 -1783
rect -275 -1817 -241 -1785
rect -275 -1887 -241 -1855
rect -275 -1889 -241 -1887
rect -275 -1955 -241 -1927
rect -275 -1961 -241 -1955
rect -275 -2023 -241 -1999
rect -275 -2033 -241 -2023
rect -275 -2091 -241 -2071
rect -275 -2105 -241 -2091
rect -275 -2159 -241 -2143
rect -275 -2177 -241 -2159
rect -275 -2227 -241 -2215
rect -275 -2249 -241 -2227
rect -275 -2295 -241 -2287
rect -275 -2321 -241 -2295
rect -275 -2363 -241 -2359
rect -275 -2393 -241 -2363
rect -275 -2465 -241 -2431
rect -17 2431 17 2465
rect -17 2363 17 2393
rect -17 2359 17 2363
rect -17 2295 17 2321
rect -17 2287 17 2295
rect -17 2227 17 2249
rect -17 2215 17 2227
rect -17 2159 17 2177
rect -17 2143 17 2159
rect -17 2091 17 2105
rect -17 2071 17 2091
rect -17 2023 17 2033
rect -17 1999 17 2023
rect -17 1955 17 1961
rect -17 1927 17 1955
rect -17 1887 17 1889
rect -17 1855 17 1887
rect -17 1785 17 1817
rect -17 1783 17 1785
rect -17 1717 17 1745
rect -17 1711 17 1717
rect -17 1649 17 1673
rect -17 1639 17 1649
rect -17 1581 17 1601
rect -17 1567 17 1581
rect -17 1513 17 1529
rect -17 1495 17 1513
rect -17 1445 17 1457
rect -17 1423 17 1445
rect -17 1377 17 1385
rect -17 1351 17 1377
rect -17 1309 17 1313
rect -17 1279 17 1309
rect -17 1207 17 1241
rect -17 1139 17 1169
rect -17 1135 17 1139
rect -17 1071 17 1097
rect -17 1063 17 1071
rect -17 1003 17 1025
rect -17 991 17 1003
rect -17 935 17 953
rect -17 919 17 935
rect -17 867 17 881
rect -17 847 17 867
rect -17 799 17 809
rect -17 775 17 799
rect -17 731 17 737
rect -17 703 17 731
rect -17 663 17 665
rect -17 631 17 663
rect -17 561 17 593
rect -17 559 17 561
rect -17 493 17 521
rect -17 487 17 493
rect -17 425 17 449
rect -17 415 17 425
rect -17 357 17 377
rect -17 343 17 357
rect -17 289 17 305
rect -17 271 17 289
rect -17 221 17 233
rect -17 199 17 221
rect -17 153 17 161
rect -17 127 17 153
rect -17 85 17 89
rect -17 55 17 85
rect -17 -17 17 17
rect -17 -85 17 -55
rect -17 -89 17 -85
rect -17 -153 17 -127
rect -17 -161 17 -153
rect -17 -221 17 -199
rect -17 -233 17 -221
rect -17 -289 17 -271
rect -17 -305 17 -289
rect -17 -357 17 -343
rect -17 -377 17 -357
rect -17 -425 17 -415
rect -17 -449 17 -425
rect -17 -493 17 -487
rect -17 -521 17 -493
rect -17 -561 17 -559
rect -17 -593 17 -561
rect -17 -663 17 -631
rect -17 -665 17 -663
rect -17 -731 17 -703
rect -17 -737 17 -731
rect -17 -799 17 -775
rect -17 -809 17 -799
rect -17 -867 17 -847
rect -17 -881 17 -867
rect -17 -935 17 -919
rect -17 -953 17 -935
rect -17 -1003 17 -991
rect -17 -1025 17 -1003
rect -17 -1071 17 -1063
rect -17 -1097 17 -1071
rect -17 -1139 17 -1135
rect -17 -1169 17 -1139
rect -17 -1241 17 -1207
rect -17 -1309 17 -1279
rect -17 -1313 17 -1309
rect -17 -1377 17 -1351
rect -17 -1385 17 -1377
rect -17 -1445 17 -1423
rect -17 -1457 17 -1445
rect -17 -1513 17 -1495
rect -17 -1529 17 -1513
rect -17 -1581 17 -1567
rect -17 -1601 17 -1581
rect -17 -1649 17 -1639
rect -17 -1673 17 -1649
rect -17 -1717 17 -1711
rect -17 -1745 17 -1717
rect -17 -1785 17 -1783
rect -17 -1817 17 -1785
rect -17 -1887 17 -1855
rect -17 -1889 17 -1887
rect -17 -1955 17 -1927
rect -17 -1961 17 -1955
rect -17 -2023 17 -1999
rect -17 -2033 17 -2023
rect -17 -2091 17 -2071
rect -17 -2105 17 -2091
rect -17 -2159 17 -2143
rect -17 -2177 17 -2159
rect -17 -2227 17 -2215
rect -17 -2249 17 -2227
rect -17 -2295 17 -2287
rect -17 -2321 17 -2295
rect -17 -2363 17 -2359
rect -17 -2393 17 -2363
rect -17 -2465 17 -2431
rect 241 2431 275 2465
rect 241 2363 275 2393
rect 241 2359 275 2363
rect 241 2295 275 2321
rect 241 2287 275 2295
rect 241 2227 275 2249
rect 241 2215 275 2227
rect 241 2159 275 2177
rect 241 2143 275 2159
rect 241 2091 275 2105
rect 241 2071 275 2091
rect 241 2023 275 2033
rect 241 1999 275 2023
rect 241 1955 275 1961
rect 241 1927 275 1955
rect 241 1887 275 1889
rect 241 1855 275 1887
rect 241 1785 275 1817
rect 241 1783 275 1785
rect 241 1717 275 1745
rect 241 1711 275 1717
rect 241 1649 275 1673
rect 241 1639 275 1649
rect 241 1581 275 1601
rect 241 1567 275 1581
rect 241 1513 275 1529
rect 241 1495 275 1513
rect 241 1445 275 1457
rect 241 1423 275 1445
rect 241 1377 275 1385
rect 241 1351 275 1377
rect 241 1309 275 1313
rect 241 1279 275 1309
rect 241 1207 275 1241
rect 241 1139 275 1169
rect 241 1135 275 1139
rect 241 1071 275 1097
rect 241 1063 275 1071
rect 241 1003 275 1025
rect 241 991 275 1003
rect 241 935 275 953
rect 241 919 275 935
rect 241 867 275 881
rect 241 847 275 867
rect 241 799 275 809
rect 241 775 275 799
rect 241 731 275 737
rect 241 703 275 731
rect 241 663 275 665
rect 241 631 275 663
rect 241 561 275 593
rect 241 559 275 561
rect 241 493 275 521
rect 241 487 275 493
rect 241 425 275 449
rect 241 415 275 425
rect 241 357 275 377
rect 241 343 275 357
rect 241 289 275 305
rect 241 271 275 289
rect 241 221 275 233
rect 241 199 275 221
rect 241 153 275 161
rect 241 127 275 153
rect 241 85 275 89
rect 241 55 275 85
rect 241 -17 275 17
rect 241 -85 275 -55
rect 241 -89 275 -85
rect 241 -153 275 -127
rect 241 -161 275 -153
rect 241 -221 275 -199
rect 241 -233 275 -221
rect 241 -289 275 -271
rect 241 -305 275 -289
rect 241 -357 275 -343
rect 241 -377 275 -357
rect 241 -425 275 -415
rect 241 -449 275 -425
rect 241 -493 275 -487
rect 241 -521 275 -493
rect 241 -561 275 -559
rect 241 -593 275 -561
rect 241 -663 275 -631
rect 241 -665 275 -663
rect 241 -731 275 -703
rect 241 -737 275 -731
rect 241 -799 275 -775
rect 241 -809 275 -799
rect 241 -867 275 -847
rect 241 -881 275 -867
rect 241 -935 275 -919
rect 241 -953 275 -935
rect 241 -1003 275 -991
rect 241 -1025 275 -1003
rect 241 -1071 275 -1063
rect 241 -1097 275 -1071
rect 241 -1139 275 -1135
rect 241 -1169 275 -1139
rect 241 -1241 275 -1207
rect 241 -1309 275 -1279
rect 241 -1313 275 -1309
rect 241 -1377 275 -1351
rect 241 -1385 275 -1377
rect 241 -1445 275 -1423
rect 241 -1457 275 -1445
rect 241 -1513 275 -1495
rect 241 -1529 275 -1513
rect 241 -1581 275 -1567
rect 241 -1601 275 -1581
rect 241 -1649 275 -1639
rect 241 -1673 275 -1649
rect 241 -1717 275 -1711
rect 241 -1745 275 -1717
rect 241 -1785 275 -1783
rect 241 -1817 275 -1785
rect 241 -1887 275 -1855
rect 241 -1889 275 -1887
rect 241 -1955 275 -1927
rect 241 -1961 275 -1955
rect 241 -2023 275 -1999
rect 241 -2033 275 -2023
rect 241 -2091 275 -2071
rect 241 -2105 275 -2091
rect 241 -2159 275 -2143
rect 241 -2177 275 -2159
rect 241 -2227 275 -2215
rect 241 -2249 275 -2227
rect 241 -2295 275 -2287
rect 241 -2321 275 -2295
rect 241 -2363 275 -2359
rect 241 -2393 275 -2363
rect 241 -2465 275 -2431
rect 499 2431 533 2465
rect 499 2363 533 2393
rect 499 2359 533 2363
rect 499 2295 533 2321
rect 499 2287 533 2295
rect 499 2227 533 2249
rect 499 2215 533 2227
rect 499 2159 533 2177
rect 499 2143 533 2159
rect 499 2091 533 2105
rect 499 2071 533 2091
rect 499 2023 533 2033
rect 499 1999 533 2023
rect 499 1955 533 1961
rect 499 1927 533 1955
rect 499 1887 533 1889
rect 499 1855 533 1887
rect 499 1785 533 1817
rect 499 1783 533 1785
rect 499 1717 533 1745
rect 499 1711 533 1717
rect 499 1649 533 1673
rect 499 1639 533 1649
rect 499 1581 533 1601
rect 499 1567 533 1581
rect 499 1513 533 1529
rect 499 1495 533 1513
rect 499 1445 533 1457
rect 499 1423 533 1445
rect 499 1377 533 1385
rect 499 1351 533 1377
rect 499 1309 533 1313
rect 499 1279 533 1309
rect 499 1207 533 1241
rect 499 1139 533 1169
rect 499 1135 533 1139
rect 499 1071 533 1097
rect 499 1063 533 1071
rect 499 1003 533 1025
rect 499 991 533 1003
rect 499 935 533 953
rect 499 919 533 935
rect 499 867 533 881
rect 499 847 533 867
rect 499 799 533 809
rect 499 775 533 799
rect 499 731 533 737
rect 499 703 533 731
rect 499 663 533 665
rect 499 631 533 663
rect 499 561 533 593
rect 499 559 533 561
rect 499 493 533 521
rect 499 487 533 493
rect 499 425 533 449
rect 499 415 533 425
rect 499 357 533 377
rect 499 343 533 357
rect 499 289 533 305
rect 499 271 533 289
rect 499 221 533 233
rect 499 199 533 221
rect 499 153 533 161
rect 499 127 533 153
rect 499 85 533 89
rect 499 55 533 85
rect 499 -17 533 17
rect 499 -85 533 -55
rect 499 -89 533 -85
rect 499 -153 533 -127
rect 499 -161 533 -153
rect 499 -221 533 -199
rect 499 -233 533 -221
rect 499 -289 533 -271
rect 499 -305 533 -289
rect 499 -357 533 -343
rect 499 -377 533 -357
rect 499 -425 533 -415
rect 499 -449 533 -425
rect 499 -493 533 -487
rect 499 -521 533 -493
rect 499 -561 533 -559
rect 499 -593 533 -561
rect 499 -663 533 -631
rect 499 -665 533 -663
rect 499 -731 533 -703
rect 499 -737 533 -731
rect 499 -799 533 -775
rect 499 -809 533 -799
rect 499 -867 533 -847
rect 499 -881 533 -867
rect 499 -935 533 -919
rect 499 -953 533 -935
rect 499 -1003 533 -991
rect 499 -1025 533 -1003
rect 499 -1071 533 -1063
rect 499 -1097 533 -1071
rect 499 -1139 533 -1135
rect 499 -1169 533 -1139
rect 499 -1241 533 -1207
rect 499 -1309 533 -1279
rect 499 -1313 533 -1309
rect 499 -1377 533 -1351
rect 499 -1385 533 -1377
rect 499 -1445 533 -1423
rect 499 -1457 533 -1445
rect 499 -1513 533 -1495
rect 499 -1529 533 -1513
rect 499 -1581 533 -1567
rect 499 -1601 533 -1581
rect 499 -1649 533 -1639
rect 499 -1673 533 -1649
rect 499 -1717 533 -1711
rect 499 -1745 533 -1717
rect 499 -1785 533 -1783
rect 499 -1817 533 -1785
rect 499 -1887 533 -1855
rect 499 -1889 533 -1887
rect 499 -1955 533 -1927
rect 499 -1961 533 -1955
rect 499 -2023 533 -1999
rect 499 -2033 533 -2023
rect 499 -2091 533 -2071
rect 499 -2105 533 -2091
rect 499 -2159 533 -2143
rect 499 -2177 533 -2159
rect 499 -2227 533 -2215
rect 499 -2249 533 -2227
rect 499 -2295 533 -2287
rect 499 -2321 533 -2295
rect 499 -2363 533 -2359
rect 499 -2393 533 -2363
rect 499 -2465 533 -2431
rect 757 2431 791 2465
rect 757 2363 791 2393
rect 757 2359 791 2363
rect 757 2295 791 2321
rect 757 2287 791 2295
rect 757 2227 791 2249
rect 757 2215 791 2227
rect 757 2159 791 2177
rect 757 2143 791 2159
rect 757 2091 791 2105
rect 757 2071 791 2091
rect 757 2023 791 2033
rect 757 1999 791 2023
rect 757 1955 791 1961
rect 757 1927 791 1955
rect 757 1887 791 1889
rect 757 1855 791 1887
rect 757 1785 791 1817
rect 757 1783 791 1785
rect 757 1717 791 1745
rect 757 1711 791 1717
rect 757 1649 791 1673
rect 757 1639 791 1649
rect 757 1581 791 1601
rect 757 1567 791 1581
rect 757 1513 791 1529
rect 757 1495 791 1513
rect 757 1445 791 1457
rect 757 1423 791 1445
rect 757 1377 791 1385
rect 757 1351 791 1377
rect 757 1309 791 1313
rect 757 1279 791 1309
rect 757 1207 791 1241
rect 757 1139 791 1169
rect 757 1135 791 1139
rect 757 1071 791 1097
rect 757 1063 791 1071
rect 757 1003 791 1025
rect 757 991 791 1003
rect 757 935 791 953
rect 757 919 791 935
rect 757 867 791 881
rect 757 847 791 867
rect 757 799 791 809
rect 757 775 791 799
rect 757 731 791 737
rect 757 703 791 731
rect 757 663 791 665
rect 757 631 791 663
rect 757 561 791 593
rect 757 559 791 561
rect 757 493 791 521
rect 757 487 791 493
rect 757 425 791 449
rect 757 415 791 425
rect 757 357 791 377
rect 757 343 791 357
rect 757 289 791 305
rect 757 271 791 289
rect 757 221 791 233
rect 757 199 791 221
rect 757 153 791 161
rect 757 127 791 153
rect 757 85 791 89
rect 757 55 791 85
rect 757 -17 791 17
rect 757 -85 791 -55
rect 757 -89 791 -85
rect 757 -153 791 -127
rect 757 -161 791 -153
rect 757 -221 791 -199
rect 757 -233 791 -221
rect 757 -289 791 -271
rect 757 -305 791 -289
rect 757 -357 791 -343
rect 757 -377 791 -357
rect 757 -425 791 -415
rect 757 -449 791 -425
rect 757 -493 791 -487
rect 757 -521 791 -493
rect 757 -561 791 -559
rect 757 -593 791 -561
rect 757 -663 791 -631
rect 757 -665 791 -663
rect 757 -731 791 -703
rect 757 -737 791 -731
rect 757 -799 791 -775
rect 757 -809 791 -799
rect 757 -867 791 -847
rect 757 -881 791 -867
rect 757 -935 791 -919
rect 757 -953 791 -935
rect 757 -1003 791 -991
rect 757 -1025 791 -1003
rect 757 -1071 791 -1063
rect 757 -1097 791 -1071
rect 757 -1139 791 -1135
rect 757 -1169 791 -1139
rect 757 -1241 791 -1207
rect 757 -1309 791 -1279
rect 757 -1313 791 -1309
rect 757 -1377 791 -1351
rect 757 -1385 791 -1377
rect 757 -1445 791 -1423
rect 757 -1457 791 -1445
rect 757 -1513 791 -1495
rect 757 -1529 791 -1513
rect 757 -1581 791 -1567
rect 757 -1601 791 -1581
rect 757 -1649 791 -1639
rect 757 -1673 791 -1649
rect 757 -1717 791 -1711
rect 757 -1745 791 -1717
rect 757 -1785 791 -1783
rect 757 -1817 791 -1785
rect 757 -1887 791 -1855
rect 757 -1889 791 -1887
rect 757 -1955 791 -1927
rect 757 -1961 791 -1955
rect 757 -2023 791 -1999
rect 757 -2033 791 -2023
rect 757 -2091 791 -2071
rect 757 -2105 791 -2091
rect 757 -2159 791 -2143
rect 757 -2177 791 -2159
rect 757 -2227 791 -2215
rect 757 -2249 791 -2227
rect 757 -2295 791 -2287
rect 757 -2321 791 -2295
rect 757 -2363 791 -2359
rect 757 -2393 791 -2363
rect 757 -2465 791 -2431
rect 1015 2431 1049 2465
rect 1015 2363 1049 2393
rect 1015 2359 1049 2363
rect 1015 2295 1049 2321
rect 1015 2287 1049 2295
rect 1015 2227 1049 2249
rect 1015 2215 1049 2227
rect 1015 2159 1049 2177
rect 1015 2143 1049 2159
rect 1015 2091 1049 2105
rect 1015 2071 1049 2091
rect 1015 2023 1049 2033
rect 1015 1999 1049 2023
rect 1015 1955 1049 1961
rect 1015 1927 1049 1955
rect 1015 1887 1049 1889
rect 1015 1855 1049 1887
rect 1015 1785 1049 1817
rect 1015 1783 1049 1785
rect 1015 1717 1049 1745
rect 1015 1711 1049 1717
rect 1015 1649 1049 1673
rect 1015 1639 1049 1649
rect 1015 1581 1049 1601
rect 1015 1567 1049 1581
rect 1015 1513 1049 1529
rect 1015 1495 1049 1513
rect 1015 1445 1049 1457
rect 1015 1423 1049 1445
rect 1015 1377 1049 1385
rect 1015 1351 1049 1377
rect 1015 1309 1049 1313
rect 1015 1279 1049 1309
rect 1015 1207 1049 1241
rect 1015 1139 1049 1169
rect 1015 1135 1049 1139
rect 1015 1071 1049 1097
rect 1015 1063 1049 1071
rect 1015 1003 1049 1025
rect 1015 991 1049 1003
rect 1015 935 1049 953
rect 1015 919 1049 935
rect 1015 867 1049 881
rect 1015 847 1049 867
rect 1015 799 1049 809
rect 1015 775 1049 799
rect 1015 731 1049 737
rect 1015 703 1049 731
rect 1015 663 1049 665
rect 1015 631 1049 663
rect 1015 561 1049 593
rect 1015 559 1049 561
rect 1015 493 1049 521
rect 1015 487 1049 493
rect 1015 425 1049 449
rect 1015 415 1049 425
rect 1015 357 1049 377
rect 1015 343 1049 357
rect 1015 289 1049 305
rect 1015 271 1049 289
rect 1015 221 1049 233
rect 1015 199 1049 221
rect 1015 153 1049 161
rect 1015 127 1049 153
rect 1015 85 1049 89
rect 1015 55 1049 85
rect 1015 -17 1049 17
rect 1015 -85 1049 -55
rect 1015 -89 1049 -85
rect 1015 -153 1049 -127
rect 1015 -161 1049 -153
rect 1015 -221 1049 -199
rect 1015 -233 1049 -221
rect 1015 -289 1049 -271
rect 1015 -305 1049 -289
rect 1015 -357 1049 -343
rect 1015 -377 1049 -357
rect 1015 -425 1049 -415
rect 1015 -449 1049 -425
rect 1015 -493 1049 -487
rect 1015 -521 1049 -493
rect 1015 -561 1049 -559
rect 1015 -593 1049 -561
rect 1015 -663 1049 -631
rect 1015 -665 1049 -663
rect 1015 -731 1049 -703
rect 1015 -737 1049 -731
rect 1015 -799 1049 -775
rect 1015 -809 1049 -799
rect 1015 -867 1049 -847
rect 1015 -881 1049 -867
rect 1015 -935 1049 -919
rect 1015 -953 1049 -935
rect 1015 -1003 1049 -991
rect 1015 -1025 1049 -1003
rect 1015 -1071 1049 -1063
rect 1015 -1097 1049 -1071
rect 1015 -1139 1049 -1135
rect 1015 -1169 1049 -1139
rect 1015 -1241 1049 -1207
rect 1015 -1309 1049 -1279
rect 1015 -1313 1049 -1309
rect 1015 -1377 1049 -1351
rect 1015 -1385 1049 -1377
rect 1015 -1445 1049 -1423
rect 1015 -1457 1049 -1445
rect 1015 -1513 1049 -1495
rect 1015 -1529 1049 -1513
rect 1015 -1581 1049 -1567
rect 1015 -1601 1049 -1581
rect 1015 -1649 1049 -1639
rect 1015 -1673 1049 -1649
rect 1015 -1717 1049 -1711
rect 1015 -1745 1049 -1717
rect 1015 -1785 1049 -1783
rect 1015 -1817 1049 -1785
rect 1015 -1887 1049 -1855
rect 1015 -1889 1049 -1887
rect 1015 -1955 1049 -1927
rect 1015 -1961 1049 -1955
rect 1015 -2023 1049 -1999
rect 1015 -2033 1049 -2023
rect 1015 -2091 1049 -2071
rect 1015 -2105 1049 -2091
rect 1015 -2159 1049 -2143
rect 1015 -2177 1049 -2159
rect 1015 -2227 1049 -2215
rect 1015 -2249 1049 -2227
rect 1015 -2295 1049 -2287
rect 1015 -2321 1049 -2295
rect 1015 -2363 1049 -2359
rect 1015 -2393 1049 -2363
rect 1015 -2465 1049 -2431
rect 1273 2431 1307 2465
rect 1273 2363 1307 2393
rect 1273 2359 1307 2363
rect 1273 2295 1307 2321
rect 1273 2287 1307 2295
rect 1273 2227 1307 2249
rect 1273 2215 1307 2227
rect 1273 2159 1307 2177
rect 1273 2143 1307 2159
rect 1273 2091 1307 2105
rect 1273 2071 1307 2091
rect 1273 2023 1307 2033
rect 1273 1999 1307 2023
rect 1273 1955 1307 1961
rect 1273 1927 1307 1955
rect 1273 1887 1307 1889
rect 1273 1855 1307 1887
rect 1273 1785 1307 1817
rect 1273 1783 1307 1785
rect 1273 1717 1307 1745
rect 1273 1711 1307 1717
rect 1273 1649 1307 1673
rect 1273 1639 1307 1649
rect 1273 1581 1307 1601
rect 1273 1567 1307 1581
rect 1273 1513 1307 1529
rect 1273 1495 1307 1513
rect 1273 1445 1307 1457
rect 1273 1423 1307 1445
rect 1273 1377 1307 1385
rect 1273 1351 1307 1377
rect 1273 1309 1307 1313
rect 1273 1279 1307 1309
rect 1273 1207 1307 1241
rect 1273 1139 1307 1169
rect 1273 1135 1307 1139
rect 1273 1071 1307 1097
rect 1273 1063 1307 1071
rect 1273 1003 1307 1025
rect 1273 991 1307 1003
rect 1273 935 1307 953
rect 1273 919 1307 935
rect 1273 867 1307 881
rect 1273 847 1307 867
rect 1273 799 1307 809
rect 1273 775 1307 799
rect 1273 731 1307 737
rect 1273 703 1307 731
rect 1273 663 1307 665
rect 1273 631 1307 663
rect 1273 561 1307 593
rect 1273 559 1307 561
rect 1273 493 1307 521
rect 1273 487 1307 493
rect 1273 425 1307 449
rect 1273 415 1307 425
rect 1273 357 1307 377
rect 1273 343 1307 357
rect 1273 289 1307 305
rect 1273 271 1307 289
rect 1273 221 1307 233
rect 1273 199 1307 221
rect 1273 153 1307 161
rect 1273 127 1307 153
rect 1273 85 1307 89
rect 1273 55 1307 85
rect 1273 -17 1307 17
rect 1273 -85 1307 -55
rect 1273 -89 1307 -85
rect 1273 -153 1307 -127
rect 1273 -161 1307 -153
rect 1273 -221 1307 -199
rect 1273 -233 1307 -221
rect 1273 -289 1307 -271
rect 1273 -305 1307 -289
rect 1273 -357 1307 -343
rect 1273 -377 1307 -357
rect 1273 -425 1307 -415
rect 1273 -449 1307 -425
rect 1273 -493 1307 -487
rect 1273 -521 1307 -493
rect 1273 -561 1307 -559
rect 1273 -593 1307 -561
rect 1273 -663 1307 -631
rect 1273 -665 1307 -663
rect 1273 -731 1307 -703
rect 1273 -737 1307 -731
rect 1273 -799 1307 -775
rect 1273 -809 1307 -799
rect 1273 -867 1307 -847
rect 1273 -881 1307 -867
rect 1273 -935 1307 -919
rect 1273 -953 1307 -935
rect 1273 -1003 1307 -991
rect 1273 -1025 1307 -1003
rect 1273 -1071 1307 -1063
rect 1273 -1097 1307 -1071
rect 1273 -1139 1307 -1135
rect 1273 -1169 1307 -1139
rect 1273 -1241 1307 -1207
rect 1273 -1309 1307 -1279
rect 1273 -1313 1307 -1309
rect 1273 -1377 1307 -1351
rect 1273 -1385 1307 -1377
rect 1273 -1445 1307 -1423
rect 1273 -1457 1307 -1445
rect 1273 -1513 1307 -1495
rect 1273 -1529 1307 -1513
rect 1273 -1581 1307 -1567
rect 1273 -1601 1307 -1581
rect 1273 -1649 1307 -1639
rect 1273 -1673 1307 -1649
rect 1273 -1717 1307 -1711
rect 1273 -1745 1307 -1717
rect 1273 -1785 1307 -1783
rect 1273 -1817 1307 -1785
rect 1273 -1887 1307 -1855
rect 1273 -1889 1307 -1887
rect 1273 -1955 1307 -1927
rect 1273 -1961 1307 -1955
rect 1273 -2023 1307 -1999
rect 1273 -2033 1307 -2023
rect 1273 -2091 1307 -2071
rect 1273 -2105 1307 -2091
rect 1273 -2159 1307 -2143
rect 1273 -2177 1307 -2159
rect 1273 -2227 1307 -2215
rect 1273 -2249 1307 -2227
rect 1273 -2295 1307 -2287
rect 1273 -2321 1307 -2295
rect 1273 -2363 1307 -2359
rect 1273 -2393 1307 -2363
rect 1273 -2465 1307 -2431
rect -1214 -2572 -1212 -2538
rect -1212 -2572 -1180 -2538
rect -1142 -2572 -1110 -2538
rect -1110 -2572 -1108 -2538
rect -956 -2572 -954 -2538
rect -954 -2572 -922 -2538
rect -884 -2572 -852 -2538
rect -852 -2572 -850 -2538
rect -698 -2572 -696 -2538
rect -696 -2572 -664 -2538
rect -626 -2572 -594 -2538
rect -594 -2572 -592 -2538
rect -440 -2572 -438 -2538
rect -438 -2572 -406 -2538
rect -368 -2572 -336 -2538
rect -336 -2572 -334 -2538
rect -182 -2572 -180 -2538
rect -180 -2572 -148 -2538
rect -110 -2572 -78 -2538
rect -78 -2572 -76 -2538
rect 76 -2572 78 -2538
rect 78 -2572 110 -2538
rect 148 -2572 180 -2538
rect 180 -2572 182 -2538
rect 334 -2572 336 -2538
rect 336 -2572 368 -2538
rect 406 -2572 438 -2538
rect 438 -2572 440 -2538
rect 592 -2572 594 -2538
rect 594 -2572 626 -2538
rect 664 -2572 696 -2538
rect 696 -2572 698 -2538
rect 850 -2572 852 -2538
rect 852 -2572 884 -2538
rect 922 -2572 954 -2538
rect 954 -2572 956 -2538
rect 1108 -2572 1110 -2538
rect 1110 -2572 1142 -2538
rect 1180 -2572 1212 -2538
rect 1212 -2572 1214 -2538
<< metal1 >>
rect -1257 2572 -1065 2578
rect -1257 2538 -1214 2572
rect -1180 2538 -1142 2572
rect -1108 2538 -1065 2572
rect -1257 2532 -1065 2538
rect -999 2572 -807 2578
rect -999 2538 -956 2572
rect -922 2538 -884 2572
rect -850 2538 -807 2572
rect -999 2532 -807 2538
rect -741 2572 -549 2578
rect -741 2538 -698 2572
rect -664 2538 -626 2572
rect -592 2538 -549 2572
rect -741 2532 -549 2538
rect -483 2572 -291 2578
rect -483 2538 -440 2572
rect -406 2538 -368 2572
rect -334 2538 -291 2572
rect -483 2532 -291 2538
rect -225 2572 -33 2578
rect -225 2538 -182 2572
rect -148 2538 -110 2572
rect -76 2538 -33 2572
rect -225 2532 -33 2538
rect 33 2572 225 2578
rect 33 2538 76 2572
rect 110 2538 148 2572
rect 182 2538 225 2572
rect 33 2532 225 2538
rect 291 2572 483 2578
rect 291 2538 334 2572
rect 368 2538 406 2572
rect 440 2538 483 2572
rect 291 2532 483 2538
rect 549 2572 741 2578
rect 549 2538 592 2572
rect 626 2538 664 2572
rect 698 2538 741 2572
rect 549 2532 741 2538
rect 807 2572 999 2578
rect 807 2538 850 2572
rect 884 2538 922 2572
rect 956 2538 999 2572
rect 807 2532 999 2538
rect 1065 2572 1257 2578
rect 1065 2538 1108 2572
rect 1142 2538 1180 2572
rect 1214 2538 1257 2572
rect 1065 2532 1257 2538
rect -1313 2465 -1267 2500
rect -1313 2431 -1307 2465
rect -1273 2431 -1267 2465
rect -1313 2393 -1267 2431
rect -1313 2359 -1307 2393
rect -1273 2359 -1267 2393
rect -1313 2321 -1267 2359
rect -1313 2287 -1307 2321
rect -1273 2287 -1267 2321
rect -1313 2249 -1267 2287
rect -1313 2215 -1307 2249
rect -1273 2215 -1267 2249
rect -1313 2177 -1267 2215
rect -1313 2143 -1307 2177
rect -1273 2143 -1267 2177
rect -1313 2105 -1267 2143
rect -1313 2071 -1307 2105
rect -1273 2071 -1267 2105
rect -1313 2033 -1267 2071
rect -1313 1999 -1307 2033
rect -1273 1999 -1267 2033
rect -1313 1961 -1267 1999
rect -1313 1927 -1307 1961
rect -1273 1927 -1267 1961
rect -1313 1889 -1267 1927
rect -1313 1855 -1307 1889
rect -1273 1855 -1267 1889
rect -1313 1817 -1267 1855
rect -1313 1783 -1307 1817
rect -1273 1783 -1267 1817
rect -1313 1745 -1267 1783
rect -1313 1711 -1307 1745
rect -1273 1711 -1267 1745
rect -1313 1673 -1267 1711
rect -1313 1639 -1307 1673
rect -1273 1639 -1267 1673
rect -1313 1601 -1267 1639
rect -1313 1567 -1307 1601
rect -1273 1567 -1267 1601
rect -1313 1529 -1267 1567
rect -1313 1495 -1307 1529
rect -1273 1495 -1267 1529
rect -1313 1457 -1267 1495
rect -1313 1423 -1307 1457
rect -1273 1423 -1267 1457
rect -1313 1385 -1267 1423
rect -1313 1351 -1307 1385
rect -1273 1351 -1267 1385
rect -1313 1313 -1267 1351
rect -1313 1279 -1307 1313
rect -1273 1279 -1267 1313
rect -1313 1241 -1267 1279
rect -1313 1207 -1307 1241
rect -1273 1207 -1267 1241
rect -1313 1169 -1267 1207
rect -1313 1135 -1307 1169
rect -1273 1135 -1267 1169
rect -1313 1097 -1267 1135
rect -1313 1063 -1307 1097
rect -1273 1063 -1267 1097
rect -1313 1025 -1267 1063
rect -1313 991 -1307 1025
rect -1273 991 -1267 1025
rect -1313 953 -1267 991
rect -1313 919 -1307 953
rect -1273 919 -1267 953
rect -1313 881 -1267 919
rect -1313 847 -1307 881
rect -1273 847 -1267 881
rect -1313 809 -1267 847
rect -1313 775 -1307 809
rect -1273 775 -1267 809
rect -1313 737 -1267 775
rect -1313 703 -1307 737
rect -1273 703 -1267 737
rect -1313 665 -1267 703
rect -1313 631 -1307 665
rect -1273 631 -1267 665
rect -1313 593 -1267 631
rect -1313 559 -1307 593
rect -1273 559 -1267 593
rect -1313 521 -1267 559
rect -1313 487 -1307 521
rect -1273 487 -1267 521
rect -1313 449 -1267 487
rect -1313 415 -1307 449
rect -1273 415 -1267 449
rect -1313 377 -1267 415
rect -1313 343 -1307 377
rect -1273 343 -1267 377
rect -1313 305 -1267 343
rect -1313 271 -1307 305
rect -1273 271 -1267 305
rect -1313 233 -1267 271
rect -1313 199 -1307 233
rect -1273 199 -1267 233
rect -1313 161 -1267 199
rect -1313 127 -1307 161
rect -1273 127 -1267 161
rect -1313 89 -1267 127
rect -1313 55 -1307 89
rect -1273 55 -1267 89
rect -1313 17 -1267 55
rect -1313 -17 -1307 17
rect -1273 -17 -1267 17
rect -1313 -55 -1267 -17
rect -1313 -89 -1307 -55
rect -1273 -89 -1267 -55
rect -1313 -127 -1267 -89
rect -1313 -161 -1307 -127
rect -1273 -161 -1267 -127
rect -1313 -199 -1267 -161
rect -1313 -233 -1307 -199
rect -1273 -233 -1267 -199
rect -1313 -271 -1267 -233
rect -1313 -305 -1307 -271
rect -1273 -305 -1267 -271
rect -1313 -343 -1267 -305
rect -1313 -377 -1307 -343
rect -1273 -377 -1267 -343
rect -1313 -415 -1267 -377
rect -1313 -449 -1307 -415
rect -1273 -449 -1267 -415
rect -1313 -487 -1267 -449
rect -1313 -521 -1307 -487
rect -1273 -521 -1267 -487
rect -1313 -559 -1267 -521
rect -1313 -593 -1307 -559
rect -1273 -593 -1267 -559
rect -1313 -631 -1267 -593
rect -1313 -665 -1307 -631
rect -1273 -665 -1267 -631
rect -1313 -703 -1267 -665
rect -1313 -737 -1307 -703
rect -1273 -737 -1267 -703
rect -1313 -775 -1267 -737
rect -1313 -809 -1307 -775
rect -1273 -809 -1267 -775
rect -1313 -847 -1267 -809
rect -1313 -881 -1307 -847
rect -1273 -881 -1267 -847
rect -1313 -919 -1267 -881
rect -1313 -953 -1307 -919
rect -1273 -953 -1267 -919
rect -1313 -991 -1267 -953
rect -1313 -1025 -1307 -991
rect -1273 -1025 -1267 -991
rect -1313 -1063 -1267 -1025
rect -1313 -1097 -1307 -1063
rect -1273 -1097 -1267 -1063
rect -1313 -1135 -1267 -1097
rect -1313 -1169 -1307 -1135
rect -1273 -1169 -1267 -1135
rect -1313 -1207 -1267 -1169
rect -1313 -1241 -1307 -1207
rect -1273 -1241 -1267 -1207
rect -1313 -1279 -1267 -1241
rect -1313 -1313 -1307 -1279
rect -1273 -1313 -1267 -1279
rect -1313 -1351 -1267 -1313
rect -1313 -1385 -1307 -1351
rect -1273 -1385 -1267 -1351
rect -1313 -1423 -1267 -1385
rect -1313 -1457 -1307 -1423
rect -1273 -1457 -1267 -1423
rect -1313 -1495 -1267 -1457
rect -1313 -1529 -1307 -1495
rect -1273 -1529 -1267 -1495
rect -1313 -1567 -1267 -1529
rect -1313 -1601 -1307 -1567
rect -1273 -1601 -1267 -1567
rect -1313 -1639 -1267 -1601
rect -1313 -1673 -1307 -1639
rect -1273 -1673 -1267 -1639
rect -1313 -1711 -1267 -1673
rect -1313 -1745 -1307 -1711
rect -1273 -1745 -1267 -1711
rect -1313 -1783 -1267 -1745
rect -1313 -1817 -1307 -1783
rect -1273 -1817 -1267 -1783
rect -1313 -1855 -1267 -1817
rect -1313 -1889 -1307 -1855
rect -1273 -1889 -1267 -1855
rect -1313 -1927 -1267 -1889
rect -1313 -1961 -1307 -1927
rect -1273 -1961 -1267 -1927
rect -1313 -1999 -1267 -1961
rect -1313 -2033 -1307 -1999
rect -1273 -2033 -1267 -1999
rect -1313 -2071 -1267 -2033
rect -1313 -2105 -1307 -2071
rect -1273 -2105 -1267 -2071
rect -1313 -2143 -1267 -2105
rect -1313 -2177 -1307 -2143
rect -1273 -2177 -1267 -2143
rect -1313 -2215 -1267 -2177
rect -1313 -2249 -1307 -2215
rect -1273 -2249 -1267 -2215
rect -1313 -2287 -1267 -2249
rect -1313 -2321 -1307 -2287
rect -1273 -2321 -1267 -2287
rect -1313 -2359 -1267 -2321
rect -1313 -2393 -1307 -2359
rect -1273 -2393 -1267 -2359
rect -1313 -2431 -1267 -2393
rect -1313 -2465 -1307 -2431
rect -1273 -2465 -1267 -2431
rect -1313 -2500 -1267 -2465
rect -1055 2465 -1009 2500
rect -1055 2431 -1049 2465
rect -1015 2431 -1009 2465
rect -1055 2393 -1009 2431
rect -1055 2359 -1049 2393
rect -1015 2359 -1009 2393
rect -1055 2321 -1009 2359
rect -1055 2287 -1049 2321
rect -1015 2287 -1009 2321
rect -1055 2249 -1009 2287
rect -1055 2215 -1049 2249
rect -1015 2215 -1009 2249
rect -1055 2177 -1009 2215
rect -1055 2143 -1049 2177
rect -1015 2143 -1009 2177
rect -1055 2105 -1009 2143
rect -1055 2071 -1049 2105
rect -1015 2071 -1009 2105
rect -1055 2033 -1009 2071
rect -1055 1999 -1049 2033
rect -1015 1999 -1009 2033
rect -1055 1961 -1009 1999
rect -1055 1927 -1049 1961
rect -1015 1927 -1009 1961
rect -1055 1889 -1009 1927
rect -1055 1855 -1049 1889
rect -1015 1855 -1009 1889
rect -1055 1817 -1009 1855
rect -1055 1783 -1049 1817
rect -1015 1783 -1009 1817
rect -1055 1745 -1009 1783
rect -1055 1711 -1049 1745
rect -1015 1711 -1009 1745
rect -1055 1673 -1009 1711
rect -1055 1639 -1049 1673
rect -1015 1639 -1009 1673
rect -1055 1601 -1009 1639
rect -1055 1567 -1049 1601
rect -1015 1567 -1009 1601
rect -1055 1529 -1009 1567
rect -1055 1495 -1049 1529
rect -1015 1495 -1009 1529
rect -1055 1457 -1009 1495
rect -1055 1423 -1049 1457
rect -1015 1423 -1009 1457
rect -1055 1385 -1009 1423
rect -1055 1351 -1049 1385
rect -1015 1351 -1009 1385
rect -1055 1313 -1009 1351
rect -1055 1279 -1049 1313
rect -1015 1279 -1009 1313
rect -1055 1241 -1009 1279
rect -1055 1207 -1049 1241
rect -1015 1207 -1009 1241
rect -1055 1169 -1009 1207
rect -1055 1135 -1049 1169
rect -1015 1135 -1009 1169
rect -1055 1097 -1009 1135
rect -1055 1063 -1049 1097
rect -1015 1063 -1009 1097
rect -1055 1025 -1009 1063
rect -1055 991 -1049 1025
rect -1015 991 -1009 1025
rect -1055 953 -1009 991
rect -1055 919 -1049 953
rect -1015 919 -1009 953
rect -1055 881 -1009 919
rect -1055 847 -1049 881
rect -1015 847 -1009 881
rect -1055 809 -1009 847
rect -1055 775 -1049 809
rect -1015 775 -1009 809
rect -1055 737 -1009 775
rect -1055 703 -1049 737
rect -1015 703 -1009 737
rect -1055 665 -1009 703
rect -1055 631 -1049 665
rect -1015 631 -1009 665
rect -1055 593 -1009 631
rect -1055 559 -1049 593
rect -1015 559 -1009 593
rect -1055 521 -1009 559
rect -1055 487 -1049 521
rect -1015 487 -1009 521
rect -1055 449 -1009 487
rect -1055 415 -1049 449
rect -1015 415 -1009 449
rect -1055 377 -1009 415
rect -1055 343 -1049 377
rect -1015 343 -1009 377
rect -1055 305 -1009 343
rect -1055 271 -1049 305
rect -1015 271 -1009 305
rect -1055 233 -1009 271
rect -1055 199 -1049 233
rect -1015 199 -1009 233
rect -1055 161 -1009 199
rect -1055 127 -1049 161
rect -1015 127 -1009 161
rect -1055 89 -1009 127
rect -1055 55 -1049 89
rect -1015 55 -1009 89
rect -1055 17 -1009 55
rect -1055 -17 -1049 17
rect -1015 -17 -1009 17
rect -1055 -55 -1009 -17
rect -1055 -89 -1049 -55
rect -1015 -89 -1009 -55
rect -1055 -127 -1009 -89
rect -1055 -161 -1049 -127
rect -1015 -161 -1009 -127
rect -1055 -199 -1009 -161
rect -1055 -233 -1049 -199
rect -1015 -233 -1009 -199
rect -1055 -271 -1009 -233
rect -1055 -305 -1049 -271
rect -1015 -305 -1009 -271
rect -1055 -343 -1009 -305
rect -1055 -377 -1049 -343
rect -1015 -377 -1009 -343
rect -1055 -415 -1009 -377
rect -1055 -449 -1049 -415
rect -1015 -449 -1009 -415
rect -1055 -487 -1009 -449
rect -1055 -521 -1049 -487
rect -1015 -521 -1009 -487
rect -1055 -559 -1009 -521
rect -1055 -593 -1049 -559
rect -1015 -593 -1009 -559
rect -1055 -631 -1009 -593
rect -1055 -665 -1049 -631
rect -1015 -665 -1009 -631
rect -1055 -703 -1009 -665
rect -1055 -737 -1049 -703
rect -1015 -737 -1009 -703
rect -1055 -775 -1009 -737
rect -1055 -809 -1049 -775
rect -1015 -809 -1009 -775
rect -1055 -847 -1009 -809
rect -1055 -881 -1049 -847
rect -1015 -881 -1009 -847
rect -1055 -919 -1009 -881
rect -1055 -953 -1049 -919
rect -1015 -953 -1009 -919
rect -1055 -991 -1009 -953
rect -1055 -1025 -1049 -991
rect -1015 -1025 -1009 -991
rect -1055 -1063 -1009 -1025
rect -1055 -1097 -1049 -1063
rect -1015 -1097 -1009 -1063
rect -1055 -1135 -1009 -1097
rect -1055 -1169 -1049 -1135
rect -1015 -1169 -1009 -1135
rect -1055 -1207 -1009 -1169
rect -1055 -1241 -1049 -1207
rect -1015 -1241 -1009 -1207
rect -1055 -1279 -1009 -1241
rect -1055 -1313 -1049 -1279
rect -1015 -1313 -1009 -1279
rect -1055 -1351 -1009 -1313
rect -1055 -1385 -1049 -1351
rect -1015 -1385 -1009 -1351
rect -1055 -1423 -1009 -1385
rect -1055 -1457 -1049 -1423
rect -1015 -1457 -1009 -1423
rect -1055 -1495 -1009 -1457
rect -1055 -1529 -1049 -1495
rect -1015 -1529 -1009 -1495
rect -1055 -1567 -1009 -1529
rect -1055 -1601 -1049 -1567
rect -1015 -1601 -1009 -1567
rect -1055 -1639 -1009 -1601
rect -1055 -1673 -1049 -1639
rect -1015 -1673 -1009 -1639
rect -1055 -1711 -1009 -1673
rect -1055 -1745 -1049 -1711
rect -1015 -1745 -1009 -1711
rect -1055 -1783 -1009 -1745
rect -1055 -1817 -1049 -1783
rect -1015 -1817 -1009 -1783
rect -1055 -1855 -1009 -1817
rect -1055 -1889 -1049 -1855
rect -1015 -1889 -1009 -1855
rect -1055 -1927 -1009 -1889
rect -1055 -1961 -1049 -1927
rect -1015 -1961 -1009 -1927
rect -1055 -1999 -1009 -1961
rect -1055 -2033 -1049 -1999
rect -1015 -2033 -1009 -1999
rect -1055 -2071 -1009 -2033
rect -1055 -2105 -1049 -2071
rect -1015 -2105 -1009 -2071
rect -1055 -2143 -1009 -2105
rect -1055 -2177 -1049 -2143
rect -1015 -2177 -1009 -2143
rect -1055 -2215 -1009 -2177
rect -1055 -2249 -1049 -2215
rect -1015 -2249 -1009 -2215
rect -1055 -2287 -1009 -2249
rect -1055 -2321 -1049 -2287
rect -1015 -2321 -1009 -2287
rect -1055 -2359 -1009 -2321
rect -1055 -2393 -1049 -2359
rect -1015 -2393 -1009 -2359
rect -1055 -2431 -1009 -2393
rect -1055 -2465 -1049 -2431
rect -1015 -2465 -1009 -2431
rect -1055 -2500 -1009 -2465
rect -797 2465 -751 2500
rect -797 2431 -791 2465
rect -757 2431 -751 2465
rect -797 2393 -751 2431
rect -797 2359 -791 2393
rect -757 2359 -751 2393
rect -797 2321 -751 2359
rect -797 2287 -791 2321
rect -757 2287 -751 2321
rect -797 2249 -751 2287
rect -797 2215 -791 2249
rect -757 2215 -751 2249
rect -797 2177 -751 2215
rect -797 2143 -791 2177
rect -757 2143 -751 2177
rect -797 2105 -751 2143
rect -797 2071 -791 2105
rect -757 2071 -751 2105
rect -797 2033 -751 2071
rect -797 1999 -791 2033
rect -757 1999 -751 2033
rect -797 1961 -751 1999
rect -797 1927 -791 1961
rect -757 1927 -751 1961
rect -797 1889 -751 1927
rect -797 1855 -791 1889
rect -757 1855 -751 1889
rect -797 1817 -751 1855
rect -797 1783 -791 1817
rect -757 1783 -751 1817
rect -797 1745 -751 1783
rect -797 1711 -791 1745
rect -757 1711 -751 1745
rect -797 1673 -751 1711
rect -797 1639 -791 1673
rect -757 1639 -751 1673
rect -797 1601 -751 1639
rect -797 1567 -791 1601
rect -757 1567 -751 1601
rect -797 1529 -751 1567
rect -797 1495 -791 1529
rect -757 1495 -751 1529
rect -797 1457 -751 1495
rect -797 1423 -791 1457
rect -757 1423 -751 1457
rect -797 1385 -751 1423
rect -797 1351 -791 1385
rect -757 1351 -751 1385
rect -797 1313 -751 1351
rect -797 1279 -791 1313
rect -757 1279 -751 1313
rect -797 1241 -751 1279
rect -797 1207 -791 1241
rect -757 1207 -751 1241
rect -797 1169 -751 1207
rect -797 1135 -791 1169
rect -757 1135 -751 1169
rect -797 1097 -751 1135
rect -797 1063 -791 1097
rect -757 1063 -751 1097
rect -797 1025 -751 1063
rect -797 991 -791 1025
rect -757 991 -751 1025
rect -797 953 -751 991
rect -797 919 -791 953
rect -757 919 -751 953
rect -797 881 -751 919
rect -797 847 -791 881
rect -757 847 -751 881
rect -797 809 -751 847
rect -797 775 -791 809
rect -757 775 -751 809
rect -797 737 -751 775
rect -797 703 -791 737
rect -757 703 -751 737
rect -797 665 -751 703
rect -797 631 -791 665
rect -757 631 -751 665
rect -797 593 -751 631
rect -797 559 -791 593
rect -757 559 -751 593
rect -797 521 -751 559
rect -797 487 -791 521
rect -757 487 -751 521
rect -797 449 -751 487
rect -797 415 -791 449
rect -757 415 -751 449
rect -797 377 -751 415
rect -797 343 -791 377
rect -757 343 -751 377
rect -797 305 -751 343
rect -797 271 -791 305
rect -757 271 -751 305
rect -797 233 -751 271
rect -797 199 -791 233
rect -757 199 -751 233
rect -797 161 -751 199
rect -797 127 -791 161
rect -757 127 -751 161
rect -797 89 -751 127
rect -797 55 -791 89
rect -757 55 -751 89
rect -797 17 -751 55
rect -797 -17 -791 17
rect -757 -17 -751 17
rect -797 -55 -751 -17
rect -797 -89 -791 -55
rect -757 -89 -751 -55
rect -797 -127 -751 -89
rect -797 -161 -791 -127
rect -757 -161 -751 -127
rect -797 -199 -751 -161
rect -797 -233 -791 -199
rect -757 -233 -751 -199
rect -797 -271 -751 -233
rect -797 -305 -791 -271
rect -757 -305 -751 -271
rect -797 -343 -751 -305
rect -797 -377 -791 -343
rect -757 -377 -751 -343
rect -797 -415 -751 -377
rect -797 -449 -791 -415
rect -757 -449 -751 -415
rect -797 -487 -751 -449
rect -797 -521 -791 -487
rect -757 -521 -751 -487
rect -797 -559 -751 -521
rect -797 -593 -791 -559
rect -757 -593 -751 -559
rect -797 -631 -751 -593
rect -797 -665 -791 -631
rect -757 -665 -751 -631
rect -797 -703 -751 -665
rect -797 -737 -791 -703
rect -757 -737 -751 -703
rect -797 -775 -751 -737
rect -797 -809 -791 -775
rect -757 -809 -751 -775
rect -797 -847 -751 -809
rect -797 -881 -791 -847
rect -757 -881 -751 -847
rect -797 -919 -751 -881
rect -797 -953 -791 -919
rect -757 -953 -751 -919
rect -797 -991 -751 -953
rect -797 -1025 -791 -991
rect -757 -1025 -751 -991
rect -797 -1063 -751 -1025
rect -797 -1097 -791 -1063
rect -757 -1097 -751 -1063
rect -797 -1135 -751 -1097
rect -797 -1169 -791 -1135
rect -757 -1169 -751 -1135
rect -797 -1207 -751 -1169
rect -797 -1241 -791 -1207
rect -757 -1241 -751 -1207
rect -797 -1279 -751 -1241
rect -797 -1313 -791 -1279
rect -757 -1313 -751 -1279
rect -797 -1351 -751 -1313
rect -797 -1385 -791 -1351
rect -757 -1385 -751 -1351
rect -797 -1423 -751 -1385
rect -797 -1457 -791 -1423
rect -757 -1457 -751 -1423
rect -797 -1495 -751 -1457
rect -797 -1529 -791 -1495
rect -757 -1529 -751 -1495
rect -797 -1567 -751 -1529
rect -797 -1601 -791 -1567
rect -757 -1601 -751 -1567
rect -797 -1639 -751 -1601
rect -797 -1673 -791 -1639
rect -757 -1673 -751 -1639
rect -797 -1711 -751 -1673
rect -797 -1745 -791 -1711
rect -757 -1745 -751 -1711
rect -797 -1783 -751 -1745
rect -797 -1817 -791 -1783
rect -757 -1817 -751 -1783
rect -797 -1855 -751 -1817
rect -797 -1889 -791 -1855
rect -757 -1889 -751 -1855
rect -797 -1927 -751 -1889
rect -797 -1961 -791 -1927
rect -757 -1961 -751 -1927
rect -797 -1999 -751 -1961
rect -797 -2033 -791 -1999
rect -757 -2033 -751 -1999
rect -797 -2071 -751 -2033
rect -797 -2105 -791 -2071
rect -757 -2105 -751 -2071
rect -797 -2143 -751 -2105
rect -797 -2177 -791 -2143
rect -757 -2177 -751 -2143
rect -797 -2215 -751 -2177
rect -797 -2249 -791 -2215
rect -757 -2249 -751 -2215
rect -797 -2287 -751 -2249
rect -797 -2321 -791 -2287
rect -757 -2321 -751 -2287
rect -797 -2359 -751 -2321
rect -797 -2393 -791 -2359
rect -757 -2393 -751 -2359
rect -797 -2431 -751 -2393
rect -797 -2465 -791 -2431
rect -757 -2465 -751 -2431
rect -797 -2500 -751 -2465
rect -539 2465 -493 2500
rect -539 2431 -533 2465
rect -499 2431 -493 2465
rect -539 2393 -493 2431
rect -539 2359 -533 2393
rect -499 2359 -493 2393
rect -539 2321 -493 2359
rect -539 2287 -533 2321
rect -499 2287 -493 2321
rect -539 2249 -493 2287
rect -539 2215 -533 2249
rect -499 2215 -493 2249
rect -539 2177 -493 2215
rect -539 2143 -533 2177
rect -499 2143 -493 2177
rect -539 2105 -493 2143
rect -539 2071 -533 2105
rect -499 2071 -493 2105
rect -539 2033 -493 2071
rect -539 1999 -533 2033
rect -499 1999 -493 2033
rect -539 1961 -493 1999
rect -539 1927 -533 1961
rect -499 1927 -493 1961
rect -539 1889 -493 1927
rect -539 1855 -533 1889
rect -499 1855 -493 1889
rect -539 1817 -493 1855
rect -539 1783 -533 1817
rect -499 1783 -493 1817
rect -539 1745 -493 1783
rect -539 1711 -533 1745
rect -499 1711 -493 1745
rect -539 1673 -493 1711
rect -539 1639 -533 1673
rect -499 1639 -493 1673
rect -539 1601 -493 1639
rect -539 1567 -533 1601
rect -499 1567 -493 1601
rect -539 1529 -493 1567
rect -539 1495 -533 1529
rect -499 1495 -493 1529
rect -539 1457 -493 1495
rect -539 1423 -533 1457
rect -499 1423 -493 1457
rect -539 1385 -493 1423
rect -539 1351 -533 1385
rect -499 1351 -493 1385
rect -539 1313 -493 1351
rect -539 1279 -533 1313
rect -499 1279 -493 1313
rect -539 1241 -493 1279
rect -539 1207 -533 1241
rect -499 1207 -493 1241
rect -539 1169 -493 1207
rect -539 1135 -533 1169
rect -499 1135 -493 1169
rect -539 1097 -493 1135
rect -539 1063 -533 1097
rect -499 1063 -493 1097
rect -539 1025 -493 1063
rect -539 991 -533 1025
rect -499 991 -493 1025
rect -539 953 -493 991
rect -539 919 -533 953
rect -499 919 -493 953
rect -539 881 -493 919
rect -539 847 -533 881
rect -499 847 -493 881
rect -539 809 -493 847
rect -539 775 -533 809
rect -499 775 -493 809
rect -539 737 -493 775
rect -539 703 -533 737
rect -499 703 -493 737
rect -539 665 -493 703
rect -539 631 -533 665
rect -499 631 -493 665
rect -539 593 -493 631
rect -539 559 -533 593
rect -499 559 -493 593
rect -539 521 -493 559
rect -539 487 -533 521
rect -499 487 -493 521
rect -539 449 -493 487
rect -539 415 -533 449
rect -499 415 -493 449
rect -539 377 -493 415
rect -539 343 -533 377
rect -499 343 -493 377
rect -539 305 -493 343
rect -539 271 -533 305
rect -499 271 -493 305
rect -539 233 -493 271
rect -539 199 -533 233
rect -499 199 -493 233
rect -539 161 -493 199
rect -539 127 -533 161
rect -499 127 -493 161
rect -539 89 -493 127
rect -539 55 -533 89
rect -499 55 -493 89
rect -539 17 -493 55
rect -539 -17 -533 17
rect -499 -17 -493 17
rect -539 -55 -493 -17
rect -539 -89 -533 -55
rect -499 -89 -493 -55
rect -539 -127 -493 -89
rect -539 -161 -533 -127
rect -499 -161 -493 -127
rect -539 -199 -493 -161
rect -539 -233 -533 -199
rect -499 -233 -493 -199
rect -539 -271 -493 -233
rect -539 -305 -533 -271
rect -499 -305 -493 -271
rect -539 -343 -493 -305
rect -539 -377 -533 -343
rect -499 -377 -493 -343
rect -539 -415 -493 -377
rect -539 -449 -533 -415
rect -499 -449 -493 -415
rect -539 -487 -493 -449
rect -539 -521 -533 -487
rect -499 -521 -493 -487
rect -539 -559 -493 -521
rect -539 -593 -533 -559
rect -499 -593 -493 -559
rect -539 -631 -493 -593
rect -539 -665 -533 -631
rect -499 -665 -493 -631
rect -539 -703 -493 -665
rect -539 -737 -533 -703
rect -499 -737 -493 -703
rect -539 -775 -493 -737
rect -539 -809 -533 -775
rect -499 -809 -493 -775
rect -539 -847 -493 -809
rect -539 -881 -533 -847
rect -499 -881 -493 -847
rect -539 -919 -493 -881
rect -539 -953 -533 -919
rect -499 -953 -493 -919
rect -539 -991 -493 -953
rect -539 -1025 -533 -991
rect -499 -1025 -493 -991
rect -539 -1063 -493 -1025
rect -539 -1097 -533 -1063
rect -499 -1097 -493 -1063
rect -539 -1135 -493 -1097
rect -539 -1169 -533 -1135
rect -499 -1169 -493 -1135
rect -539 -1207 -493 -1169
rect -539 -1241 -533 -1207
rect -499 -1241 -493 -1207
rect -539 -1279 -493 -1241
rect -539 -1313 -533 -1279
rect -499 -1313 -493 -1279
rect -539 -1351 -493 -1313
rect -539 -1385 -533 -1351
rect -499 -1385 -493 -1351
rect -539 -1423 -493 -1385
rect -539 -1457 -533 -1423
rect -499 -1457 -493 -1423
rect -539 -1495 -493 -1457
rect -539 -1529 -533 -1495
rect -499 -1529 -493 -1495
rect -539 -1567 -493 -1529
rect -539 -1601 -533 -1567
rect -499 -1601 -493 -1567
rect -539 -1639 -493 -1601
rect -539 -1673 -533 -1639
rect -499 -1673 -493 -1639
rect -539 -1711 -493 -1673
rect -539 -1745 -533 -1711
rect -499 -1745 -493 -1711
rect -539 -1783 -493 -1745
rect -539 -1817 -533 -1783
rect -499 -1817 -493 -1783
rect -539 -1855 -493 -1817
rect -539 -1889 -533 -1855
rect -499 -1889 -493 -1855
rect -539 -1927 -493 -1889
rect -539 -1961 -533 -1927
rect -499 -1961 -493 -1927
rect -539 -1999 -493 -1961
rect -539 -2033 -533 -1999
rect -499 -2033 -493 -1999
rect -539 -2071 -493 -2033
rect -539 -2105 -533 -2071
rect -499 -2105 -493 -2071
rect -539 -2143 -493 -2105
rect -539 -2177 -533 -2143
rect -499 -2177 -493 -2143
rect -539 -2215 -493 -2177
rect -539 -2249 -533 -2215
rect -499 -2249 -493 -2215
rect -539 -2287 -493 -2249
rect -539 -2321 -533 -2287
rect -499 -2321 -493 -2287
rect -539 -2359 -493 -2321
rect -539 -2393 -533 -2359
rect -499 -2393 -493 -2359
rect -539 -2431 -493 -2393
rect -539 -2465 -533 -2431
rect -499 -2465 -493 -2431
rect -539 -2500 -493 -2465
rect -281 2465 -235 2500
rect -281 2431 -275 2465
rect -241 2431 -235 2465
rect -281 2393 -235 2431
rect -281 2359 -275 2393
rect -241 2359 -235 2393
rect -281 2321 -235 2359
rect -281 2287 -275 2321
rect -241 2287 -235 2321
rect -281 2249 -235 2287
rect -281 2215 -275 2249
rect -241 2215 -235 2249
rect -281 2177 -235 2215
rect -281 2143 -275 2177
rect -241 2143 -235 2177
rect -281 2105 -235 2143
rect -281 2071 -275 2105
rect -241 2071 -235 2105
rect -281 2033 -235 2071
rect -281 1999 -275 2033
rect -241 1999 -235 2033
rect -281 1961 -235 1999
rect -281 1927 -275 1961
rect -241 1927 -235 1961
rect -281 1889 -235 1927
rect -281 1855 -275 1889
rect -241 1855 -235 1889
rect -281 1817 -235 1855
rect -281 1783 -275 1817
rect -241 1783 -235 1817
rect -281 1745 -235 1783
rect -281 1711 -275 1745
rect -241 1711 -235 1745
rect -281 1673 -235 1711
rect -281 1639 -275 1673
rect -241 1639 -235 1673
rect -281 1601 -235 1639
rect -281 1567 -275 1601
rect -241 1567 -235 1601
rect -281 1529 -235 1567
rect -281 1495 -275 1529
rect -241 1495 -235 1529
rect -281 1457 -235 1495
rect -281 1423 -275 1457
rect -241 1423 -235 1457
rect -281 1385 -235 1423
rect -281 1351 -275 1385
rect -241 1351 -235 1385
rect -281 1313 -235 1351
rect -281 1279 -275 1313
rect -241 1279 -235 1313
rect -281 1241 -235 1279
rect -281 1207 -275 1241
rect -241 1207 -235 1241
rect -281 1169 -235 1207
rect -281 1135 -275 1169
rect -241 1135 -235 1169
rect -281 1097 -235 1135
rect -281 1063 -275 1097
rect -241 1063 -235 1097
rect -281 1025 -235 1063
rect -281 991 -275 1025
rect -241 991 -235 1025
rect -281 953 -235 991
rect -281 919 -275 953
rect -241 919 -235 953
rect -281 881 -235 919
rect -281 847 -275 881
rect -241 847 -235 881
rect -281 809 -235 847
rect -281 775 -275 809
rect -241 775 -235 809
rect -281 737 -235 775
rect -281 703 -275 737
rect -241 703 -235 737
rect -281 665 -235 703
rect -281 631 -275 665
rect -241 631 -235 665
rect -281 593 -235 631
rect -281 559 -275 593
rect -241 559 -235 593
rect -281 521 -235 559
rect -281 487 -275 521
rect -241 487 -235 521
rect -281 449 -235 487
rect -281 415 -275 449
rect -241 415 -235 449
rect -281 377 -235 415
rect -281 343 -275 377
rect -241 343 -235 377
rect -281 305 -235 343
rect -281 271 -275 305
rect -241 271 -235 305
rect -281 233 -235 271
rect -281 199 -275 233
rect -241 199 -235 233
rect -281 161 -235 199
rect -281 127 -275 161
rect -241 127 -235 161
rect -281 89 -235 127
rect -281 55 -275 89
rect -241 55 -235 89
rect -281 17 -235 55
rect -281 -17 -275 17
rect -241 -17 -235 17
rect -281 -55 -235 -17
rect -281 -89 -275 -55
rect -241 -89 -235 -55
rect -281 -127 -235 -89
rect -281 -161 -275 -127
rect -241 -161 -235 -127
rect -281 -199 -235 -161
rect -281 -233 -275 -199
rect -241 -233 -235 -199
rect -281 -271 -235 -233
rect -281 -305 -275 -271
rect -241 -305 -235 -271
rect -281 -343 -235 -305
rect -281 -377 -275 -343
rect -241 -377 -235 -343
rect -281 -415 -235 -377
rect -281 -449 -275 -415
rect -241 -449 -235 -415
rect -281 -487 -235 -449
rect -281 -521 -275 -487
rect -241 -521 -235 -487
rect -281 -559 -235 -521
rect -281 -593 -275 -559
rect -241 -593 -235 -559
rect -281 -631 -235 -593
rect -281 -665 -275 -631
rect -241 -665 -235 -631
rect -281 -703 -235 -665
rect -281 -737 -275 -703
rect -241 -737 -235 -703
rect -281 -775 -235 -737
rect -281 -809 -275 -775
rect -241 -809 -235 -775
rect -281 -847 -235 -809
rect -281 -881 -275 -847
rect -241 -881 -235 -847
rect -281 -919 -235 -881
rect -281 -953 -275 -919
rect -241 -953 -235 -919
rect -281 -991 -235 -953
rect -281 -1025 -275 -991
rect -241 -1025 -235 -991
rect -281 -1063 -235 -1025
rect -281 -1097 -275 -1063
rect -241 -1097 -235 -1063
rect -281 -1135 -235 -1097
rect -281 -1169 -275 -1135
rect -241 -1169 -235 -1135
rect -281 -1207 -235 -1169
rect -281 -1241 -275 -1207
rect -241 -1241 -235 -1207
rect -281 -1279 -235 -1241
rect -281 -1313 -275 -1279
rect -241 -1313 -235 -1279
rect -281 -1351 -235 -1313
rect -281 -1385 -275 -1351
rect -241 -1385 -235 -1351
rect -281 -1423 -235 -1385
rect -281 -1457 -275 -1423
rect -241 -1457 -235 -1423
rect -281 -1495 -235 -1457
rect -281 -1529 -275 -1495
rect -241 -1529 -235 -1495
rect -281 -1567 -235 -1529
rect -281 -1601 -275 -1567
rect -241 -1601 -235 -1567
rect -281 -1639 -235 -1601
rect -281 -1673 -275 -1639
rect -241 -1673 -235 -1639
rect -281 -1711 -235 -1673
rect -281 -1745 -275 -1711
rect -241 -1745 -235 -1711
rect -281 -1783 -235 -1745
rect -281 -1817 -275 -1783
rect -241 -1817 -235 -1783
rect -281 -1855 -235 -1817
rect -281 -1889 -275 -1855
rect -241 -1889 -235 -1855
rect -281 -1927 -235 -1889
rect -281 -1961 -275 -1927
rect -241 -1961 -235 -1927
rect -281 -1999 -235 -1961
rect -281 -2033 -275 -1999
rect -241 -2033 -235 -1999
rect -281 -2071 -235 -2033
rect -281 -2105 -275 -2071
rect -241 -2105 -235 -2071
rect -281 -2143 -235 -2105
rect -281 -2177 -275 -2143
rect -241 -2177 -235 -2143
rect -281 -2215 -235 -2177
rect -281 -2249 -275 -2215
rect -241 -2249 -235 -2215
rect -281 -2287 -235 -2249
rect -281 -2321 -275 -2287
rect -241 -2321 -235 -2287
rect -281 -2359 -235 -2321
rect -281 -2393 -275 -2359
rect -241 -2393 -235 -2359
rect -281 -2431 -235 -2393
rect -281 -2465 -275 -2431
rect -241 -2465 -235 -2431
rect -281 -2500 -235 -2465
rect -23 2465 23 2500
rect -23 2431 -17 2465
rect 17 2431 23 2465
rect -23 2393 23 2431
rect -23 2359 -17 2393
rect 17 2359 23 2393
rect -23 2321 23 2359
rect -23 2287 -17 2321
rect 17 2287 23 2321
rect -23 2249 23 2287
rect -23 2215 -17 2249
rect 17 2215 23 2249
rect -23 2177 23 2215
rect -23 2143 -17 2177
rect 17 2143 23 2177
rect -23 2105 23 2143
rect -23 2071 -17 2105
rect 17 2071 23 2105
rect -23 2033 23 2071
rect -23 1999 -17 2033
rect 17 1999 23 2033
rect -23 1961 23 1999
rect -23 1927 -17 1961
rect 17 1927 23 1961
rect -23 1889 23 1927
rect -23 1855 -17 1889
rect 17 1855 23 1889
rect -23 1817 23 1855
rect -23 1783 -17 1817
rect 17 1783 23 1817
rect -23 1745 23 1783
rect -23 1711 -17 1745
rect 17 1711 23 1745
rect -23 1673 23 1711
rect -23 1639 -17 1673
rect 17 1639 23 1673
rect -23 1601 23 1639
rect -23 1567 -17 1601
rect 17 1567 23 1601
rect -23 1529 23 1567
rect -23 1495 -17 1529
rect 17 1495 23 1529
rect -23 1457 23 1495
rect -23 1423 -17 1457
rect 17 1423 23 1457
rect -23 1385 23 1423
rect -23 1351 -17 1385
rect 17 1351 23 1385
rect -23 1313 23 1351
rect -23 1279 -17 1313
rect 17 1279 23 1313
rect -23 1241 23 1279
rect -23 1207 -17 1241
rect 17 1207 23 1241
rect -23 1169 23 1207
rect -23 1135 -17 1169
rect 17 1135 23 1169
rect -23 1097 23 1135
rect -23 1063 -17 1097
rect 17 1063 23 1097
rect -23 1025 23 1063
rect -23 991 -17 1025
rect 17 991 23 1025
rect -23 953 23 991
rect -23 919 -17 953
rect 17 919 23 953
rect -23 881 23 919
rect -23 847 -17 881
rect 17 847 23 881
rect -23 809 23 847
rect -23 775 -17 809
rect 17 775 23 809
rect -23 737 23 775
rect -23 703 -17 737
rect 17 703 23 737
rect -23 665 23 703
rect -23 631 -17 665
rect 17 631 23 665
rect -23 593 23 631
rect -23 559 -17 593
rect 17 559 23 593
rect -23 521 23 559
rect -23 487 -17 521
rect 17 487 23 521
rect -23 449 23 487
rect -23 415 -17 449
rect 17 415 23 449
rect -23 377 23 415
rect -23 343 -17 377
rect 17 343 23 377
rect -23 305 23 343
rect -23 271 -17 305
rect 17 271 23 305
rect -23 233 23 271
rect -23 199 -17 233
rect 17 199 23 233
rect -23 161 23 199
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -199 23 -161
rect -23 -233 -17 -199
rect 17 -233 23 -199
rect -23 -271 23 -233
rect -23 -305 -17 -271
rect 17 -305 23 -271
rect -23 -343 23 -305
rect -23 -377 -17 -343
rect 17 -377 23 -343
rect -23 -415 23 -377
rect -23 -449 -17 -415
rect 17 -449 23 -415
rect -23 -487 23 -449
rect -23 -521 -17 -487
rect 17 -521 23 -487
rect -23 -559 23 -521
rect -23 -593 -17 -559
rect 17 -593 23 -559
rect -23 -631 23 -593
rect -23 -665 -17 -631
rect 17 -665 23 -631
rect -23 -703 23 -665
rect -23 -737 -17 -703
rect 17 -737 23 -703
rect -23 -775 23 -737
rect -23 -809 -17 -775
rect 17 -809 23 -775
rect -23 -847 23 -809
rect -23 -881 -17 -847
rect 17 -881 23 -847
rect -23 -919 23 -881
rect -23 -953 -17 -919
rect 17 -953 23 -919
rect -23 -991 23 -953
rect -23 -1025 -17 -991
rect 17 -1025 23 -991
rect -23 -1063 23 -1025
rect -23 -1097 -17 -1063
rect 17 -1097 23 -1063
rect -23 -1135 23 -1097
rect -23 -1169 -17 -1135
rect 17 -1169 23 -1135
rect -23 -1207 23 -1169
rect -23 -1241 -17 -1207
rect 17 -1241 23 -1207
rect -23 -1279 23 -1241
rect -23 -1313 -17 -1279
rect 17 -1313 23 -1279
rect -23 -1351 23 -1313
rect -23 -1385 -17 -1351
rect 17 -1385 23 -1351
rect -23 -1423 23 -1385
rect -23 -1457 -17 -1423
rect 17 -1457 23 -1423
rect -23 -1495 23 -1457
rect -23 -1529 -17 -1495
rect 17 -1529 23 -1495
rect -23 -1567 23 -1529
rect -23 -1601 -17 -1567
rect 17 -1601 23 -1567
rect -23 -1639 23 -1601
rect -23 -1673 -17 -1639
rect 17 -1673 23 -1639
rect -23 -1711 23 -1673
rect -23 -1745 -17 -1711
rect 17 -1745 23 -1711
rect -23 -1783 23 -1745
rect -23 -1817 -17 -1783
rect 17 -1817 23 -1783
rect -23 -1855 23 -1817
rect -23 -1889 -17 -1855
rect 17 -1889 23 -1855
rect -23 -1927 23 -1889
rect -23 -1961 -17 -1927
rect 17 -1961 23 -1927
rect -23 -1999 23 -1961
rect -23 -2033 -17 -1999
rect 17 -2033 23 -1999
rect -23 -2071 23 -2033
rect -23 -2105 -17 -2071
rect 17 -2105 23 -2071
rect -23 -2143 23 -2105
rect -23 -2177 -17 -2143
rect 17 -2177 23 -2143
rect -23 -2215 23 -2177
rect -23 -2249 -17 -2215
rect 17 -2249 23 -2215
rect -23 -2287 23 -2249
rect -23 -2321 -17 -2287
rect 17 -2321 23 -2287
rect -23 -2359 23 -2321
rect -23 -2393 -17 -2359
rect 17 -2393 23 -2359
rect -23 -2431 23 -2393
rect -23 -2465 -17 -2431
rect 17 -2465 23 -2431
rect -23 -2500 23 -2465
rect 235 2465 281 2500
rect 235 2431 241 2465
rect 275 2431 281 2465
rect 235 2393 281 2431
rect 235 2359 241 2393
rect 275 2359 281 2393
rect 235 2321 281 2359
rect 235 2287 241 2321
rect 275 2287 281 2321
rect 235 2249 281 2287
rect 235 2215 241 2249
rect 275 2215 281 2249
rect 235 2177 281 2215
rect 235 2143 241 2177
rect 275 2143 281 2177
rect 235 2105 281 2143
rect 235 2071 241 2105
rect 275 2071 281 2105
rect 235 2033 281 2071
rect 235 1999 241 2033
rect 275 1999 281 2033
rect 235 1961 281 1999
rect 235 1927 241 1961
rect 275 1927 281 1961
rect 235 1889 281 1927
rect 235 1855 241 1889
rect 275 1855 281 1889
rect 235 1817 281 1855
rect 235 1783 241 1817
rect 275 1783 281 1817
rect 235 1745 281 1783
rect 235 1711 241 1745
rect 275 1711 281 1745
rect 235 1673 281 1711
rect 235 1639 241 1673
rect 275 1639 281 1673
rect 235 1601 281 1639
rect 235 1567 241 1601
rect 275 1567 281 1601
rect 235 1529 281 1567
rect 235 1495 241 1529
rect 275 1495 281 1529
rect 235 1457 281 1495
rect 235 1423 241 1457
rect 275 1423 281 1457
rect 235 1385 281 1423
rect 235 1351 241 1385
rect 275 1351 281 1385
rect 235 1313 281 1351
rect 235 1279 241 1313
rect 275 1279 281 1313
rect 235 1241 281 1279
rect 235 1207 241 1241
rect 275 1207 281 1241
rect 235 1169 281 1207
rect 235 1135 241 1169
rect 275 1135 281 1169
rect 235 1097 281 1135
rect 235 1063 241 1097
rect 275 1063 281 1097
rect 235 1025 281 1063
rect 235 991 241 1025
rect 275 991 281 1025
rect 235 953 281 991
rect 235 919 241 953
rect 275 919 281 953
rect 235 881 281 919
rect 235 847 241 881
rect 275 847 281 881
rect 235 809 281 847
rect 235 775 241 809
rect 275 775 281 809
rect 235 737 281 775
rect 235 703 241 737
rect 275 703 281 737
rect 235 665 281 703
rect 235 631 241 665
rect 275 631 281 665
rect 235 593 281 631
rect 235 559 241 593
rect 275 559 281 593
rect 235 521 281 559
rect 235 487 241 521
rect 275 487 281 521
rect 235 449 281 487
rect 235 415 241 449
rect 275 415 281 449
rect 235 377 281 415
rect 235 343 241 377
rect 275 343 281 377
rect 235 305 281 343
rect 235 271 241 305
rect 275 271 281 305
rect 235 233 281 271
rect 235 199 241 233
rect 275 199 281 233
rect 235 161 281 199
rect 235 127 241 161
rect 275 127 281 161
rect 235 89 281 127
rect 235 55 241 89
rect 275 55 281 89
rect 235 17 281 55
rect 235 -17 241 17
rect 275 -17 281 17
rect 235 -55 281 -17
rect 235 -89 241 -55
rect 275 -89 281 -55
rect 235 -127 281 -89
rect 235 -161 241 -127
rect 275 -161 281 -127
rect 235 -199 281 -161
rect 235 -233 241 -199
rect 275 -233 281 -199
rect 235 -271 281 -233
rect 235 -305 241 -271
rect 275 -305 281 -271
rect 235 -343 281 -305
rect 235 -377 241 -343
rect 275 -377 281 -343
rect 235 -415 281 -377
rect 235 -449 241 -415
rect 275 -449 281 -415
rect 235 -487 281 -449
rect 235 -521 241 -487
rect 275 -521 281 -487
rect 235 -559 281 -521
rect 235 -593 241 -559
rect 275 -593 281 -559
rect 235 -631 281 -593
rect 235 -665 241 -631
rect 275 -665 281 -631
rect 235 -703 281 -665
rect 235 -737 241 -703
rect 275 -737 281 -703
rect 235 -775 281 -737
rect 235 -809 241 -775
rect 275 -809 281 -775
rect 235 -847 281 -809
rect 235 -881 241 -847
rect 275 -881 281 -847
rect 235 -919 281 -881
rect 235 -953 241 -919
rect 275 -953 281 -919
rect 235 -991 281 -953
rect 235 -1025 241 -991
rect 275 -1025 281 -991
rect 235 -1063 281 -1025
rect 235 -1097 241 -1063
rect 275 -1097 281 -1063
rect 235 -1135 281 -1097
rect 235 -1169 241 -1135
rect 275 -1169 281 -1135
rect 235 -1207 281 -1169
rect 235 -1241 241 -1207
rect 275 -1241 281 -1207
rect 235 -1279 281 -1241
rect 235 -1313 241 -1279
rect 275 -1313 281 -1279
rect 235 -1351 281 -1313
rect 235 -1385 241 -1351
rect 275 -1385 281 -1351
rect 235 -1423 281 -1385
rect 235 -1457 241 -1423
rect 275 -1457 281 -1423
rect 235 -1495 281 -1457
rect 235 -1529 241 -1495
rect 275 -1529 281 -1495
rect 235 -1567 281 -1529
rect 235 -1601 241 -1567
rect 275 -1601 281 -1567
rect 235 -1639 281 -1601
rect 235 -1673 241 -1639
rect 275 -1673 281 -1639
rect 235 -1711 281 -1673
rect 235 -1745 241 -1711
rect 275 -1745 281 -1711
rect 235 -1783 281 -1745
rect 235 -1817 241 -1783
rect 275 -1817 281 -1783
rect 235 -1855 281 -1817
rect 235 -1889 241 -1855
rect 275 -1889 281 -1855
rect 235 -1927 281 -1889
rect 235 -1961 241 -1927
rect 275 -1961 281 -1927
rect 235 -1999 281 -1961
rect 235 -2033 241 -1999
rect 275 -2033 281 -1999
rect 235 -2071 281 -2033
rect 235 -2105 241 -2071
rect 275 -2105 281 -2071
rect 235 -2143 281 -2105
rect 235 -2177 241 -2143
rect 275 -2177 281 -2143
rect 235 -2215 281 -2177
rect 235 -2249 241 -2215
rect 275 -2249 281 -2215
rect 235 -2287 281 -2249
rect 235 -2321 241 -2287
rect 275 -2321 281 -2287
rect 235 -2359 281 -2321
rect 235 -2393 241 -2359
rect 275 -2393 281 -2359
rect 235 -2431 281 -2393
rect 235 -2465 241 -2431
rect 275 -2465 281 -2431
rect 235 -2500 281 -2465
rect 493 2465 539 2500
rect 493 2431 499 2465
rect 533 2431 539 2465
rect 493 2393 539 2431
rect 493 2359 499 2393
rect 533 2359 539 2393
rect 493 2321 539 2359
rect 493 2287 499 2321
rect 533 2287 539 2321
rect 493 2249 539 2287
rect 493 2215 499 2249
rect 533 2215 539 2249
rect 493 2177 539 2215
rect 493 2143 499 2177
rect 533 2143 539 2177
rect 493 2105 539 2143
rect 493 2071 499 2105
rect 533 2071 539 2105
rect 493 2033 539 2071
rect 493 1999 499 2033
rect 533 1999 539 2033
rect 493 1961 539 1999
rect 493 1927 499 1961
rect 533 1927 539 1961
rect 493 1889 539 1927
rect 493 1855 499 1889
rect 533 1855 539 1889
rect 493 1817 539 1855
rect 493 1783 499 1817
rect 533 1783 539 1817
rect 493 1745 539 1783
rect 493 1711 499 1745
rect 533 1711 539 1745
rect 493 1673 539 1711
rect 493 1639 499 1673
rect 533 1639 539 1673
rect 493 1601 539 1639
rect 493 1567 499 1601
rect 533 1567 539 1601
rect 493 1529 539 1567
rect 493 1495 499 1529
rect 533 1495 539 1529
rect 493 1457 539 1495
rect 493 1423 499 1457
rect 533 1423 539 1457
rect 493 1385 539 1423
rect 493 1351 499 1385
rect 533 1351 539 1385
rect 493 1313 539 1351
rect 493 1279 499 1313
rect 533 1279 539 1313
rect 493 1241 539 1279
rect 493 1207 499 1241
rect 533 1207 539 1241
rect 493 1169 539 1207
rect 493 1135 499 1169
rect 533 1135 539 1169
rect 493 1097 539 1135
rect 493 1063 499 1097
rect 533 1063 539 1097
rect 493 1025 539 1063
rect 493 991 499 1025
rect 533 991 539 1025
rect 493 953 539 991
rect 493 919 499 953
rect 533 919 539 953
rect 493 881 539 919
rect 493 847 499 881
rect 533 847 539 881
rect 493 809 539 847
rect 493 775 499 809
rect 533 775 539 809
rect 493 737 539 775
rect 493 703 499 737
rect 533 703 539 737
rect 493 665 539 703
rect 493 631 499 665
rect 533 631 539 665
rect 493 593 539 631
rect 493 559 499 593
rect 533 559 539 593
rect 493 521 539 559
rect 493 487 499 521
rect 533 487 539 521
rect 493 449 539 487
rect 493 415 499 449
rect 533 415 539 449
rect 493 377 539 415
rect 493 343 499 377
rect 533 343 539 377
rect 493 305 539 343
rect 493 271 499 305
rect 533 271 539 305
rect 493 233 539 271
rect 493 199 499 233
rect 533 199 539 233
rect 493 161 539 199
rect 493 127 499 161
rect 533 127 539 161
rect 493 89 539 127
rect 493 55 499 89
rect 533 55 539 89
rect 493 17 539 55
rect 493 -17 499 17
rect 533 -17 539 17
rect 493 -55 539 -17
rect 493 -89 499 -55
rect 533 -89 539 -55
rect 493 -127 539 -89
rect 493 -161 499 -127
rect 533 -161 539 -127
rect 493 -199 539 -161
rect 493 -233 499 -199
rect 533 -233 539 -199
rect 493 -271 539 -233
rect 493 -305 499 -271
rect 533 -305 539 -271
rect 493 -343 539 -305
rect 493 -377 499 -343
rect 533 -377 539 -343
rect 493 -415 539 -377
rect 493 -449 499 -415
rect 533 -449 539 -415
rect 493 -487 539 -449
rect 493 -521 499 -487
rect 533 -521 539 -487
rect 493 -559 539 -521
rect 493 -593 499 -559
rect 533 -593 539 -559
rect 493 -631 539 -593
rect 493 -665 499 -631
rect 533 -665 539 -631
rect 493 -703 539 -665
rect 493 -737 499 -703
rect 533 -737 539 -703
rect 493 -775 539 -737
rect 493 -809 499 -775
rect 533 -809 539 -775
rect 493 -847 539 -809
rect 493 -881 499 -847
rect 533 -881 539 -847
rect 493 -919 539 -881
rect 493 -953 499 -919
rect 533 -953 539 -919
rect 493 -991 539 -953
rect 493 -1025 499 -991
rect 533 -1025 539 -991
rect 493 -1063 539 -1025
rect 493 -1097 499 -1063
rect 533 -1097 539 -1063
rect 493 -1135 539 -1097
rect 493 -1169 499 -1135
rect 533 -1169 539 -1135
rect 493 -1207 539 -1169
rect 493 -1241 499 -1207
rect 533 -1241 539 -1207
rect 493 -1279 539 -1241
rect 493 -1313 499 -1279
rect 533 -1313 539 -1279
rect 493 -1351 539 -1313
rect 493 -1385 499 -1351
rect 533 -1385 539 -1351
rect 493 -1423 539 -1385
rect 493 -1457 499 -1423
rect 533 -1457 539 -1423
rect 493 -1495 539 -1457
rect 493 -1529 499 -1495
rect 533 -1529 539 -1495
rect 493 -1567 539 -1529
rect 493 -1601 499 -1567
rect 533 -1601 539 -1567
rect 493 -1639 539 -1601
rect 493 -1673 499 -1639
rect 533 -1673 539 -1639
rect 493 -1711 539 -1673
rect 493 -1745 499 -1711
rect 533 -1745 539 -1711
rect 493 -1783 539 -1745
rect 493 -1817 499 -1783
rect 533 -1817 539 -1783
rect 493 -1855 539 -1817
rect 493 -1889 499 -1855
rect 533 -1889 539 -1855
rect 493 -1927 539 -1889
rect 493 -1961 499 -1927
rect 533 -1961 539 -1927
rect 493 -1999 539 -1961
rect 493 -2033 499 -1999
rect 533 -2033 539 -1999
rect 493 -2071 539 -2033
rect 493 -2105 499 -2071
rect 533 -2105 539 -2071
rect 493 -2143 539 -2105
rect 493 -2177 499 -2143
rect 533 -2177 539 -2143
rect 493 -2215 539 -2177
rect 493 -2249 499 -2215
rect 533 -2249 539 -2215
rect 493 -2287 539 -2249
rect 493 -2321 499 -2287
rect 533 -2321 539 -2287
rect 493 -2359 539 -2321
rect 493 -2393 499 -2359
rect 533 -2393 539 -2359
rect 493 -2431 539 -2393
rect 493 -2465 499 -2431
rect 533 -2465 539 -2431
rect 493 -2500 539 -2465
rect 751 2465 797 2500
rect 751 2431 757 2465
rect 791 2431 797 2465
rect 751 2393 797 2431
rect 751 2359 757 2393
rect 791 2359 797 2393
rect 751 2321 797 2359
rect 751 2287 757 2321
rect 791 2287 797 2321
rect 751 2249 797 2287
rect 751 2215 757 2249
rect 791 2215 797 2249
rect 751 2177 797 2215
rect 751 2143 757 2177
rect 791 2143 797 2177
rect 751 2105 797 2143
rect 751 2071 757 2105
rect 791 2071 797 2105
rect 751 2033 797 2071
rect 751 1999 757 2033
rect 791 1999 797 2033
rect 751 1961 797 1999
rect 751 1927 757 1961
rect 791 1927 797 1961
rect 751 1889 797 1927
rect 751 1855 757 1889
rect 791 1855 797 1889
rect 751 1817 797 1855
rect 751 1783 757 1817
rect 791 1783 797 1817
rect 751 1745 797 1783
rect 751 1711 757 1745
rect 791 1711 797 1745
rect 751 1673 797 1711
rect 751 1639 757 1673
rect 791 1639 797 1673
rect 751 1601 797 1639
rect 751 1567 757 1601
rect 791 1567 797 1601
rect 751 1529 797 1567
rect 751 1495 757 1529
rect 791 1495 797 1529
rect 751 1457 797 1495
rect 751 1423 757 1457
rect 791 1423 797 1457
rect 751 1385 797 1423
rect 751 1351 757 1385
rect 791 1351 797 1385
rect 751 1313 797 1351
rect 751 1279 757 1313
rect 791 1279 797 1313
rect 751 1241 797 1279
rect 751 1207 757 1241
rect 791 1207 797 1241
rect 751 1169 797 1207
rect 751 1135 757 1169
rect 791 1135 797 1169
rect 751 1097 797 1135
rect 751 1063 757 1097
rect 791 1063 797 1097
rect 751 1025 797 1063
rect 751 991 757 1025
rect 791 991 797 1025
rect 751 953 797 991
rect 751 919 757 953
rect 791 919 797 953
rect 751 881 797 919
rect 751 847 757 881
rect 791 847 797 881
rect 751 809 797 847
rect 751 775 757 809
rect 791 775 797 809
rect 751 737 797 775
rect 751 703 757 737
rect 791 703 797 737
rect 751 665 797 703
rect 751 631 757 665
rect 791 631 797 665
rect 751 593 797 631
rect 751 559 757 593
rect 791 559 797 593
rect 751 521 797 559
rect 751 487 757 521
rect 791 487 797 521
rect 751 449 797 487
rect 751 415 757 449
rect 791 415 797 449
rect 751 377 797 415
rect 751 343 757 377
rect 791 343 797 377
rect 751 305 797 343
rect 751 271 757 305
rect 791 271 797 305
rect 751 233 797 271
rect 751 199 757 233
rect 791 199 797 233
rect 751 161 797 199
rect 751 127 757 161
rect 791 127 797 161
rect 751 89 797 127
rect 751 55 757 89
rect 791 55 797 89
rect 751 17 797 55
rect 751 -17 757 17
rect 791 -17 797 17
rect 751 -55 797 -17
rect 751 -89 757 -55
rect 791 -89 797 -55
rect 751 -127 797 -89
rect 751 -161 757 -127
rect 791 -161 797 -127
rect 751 -199 797 -161
rect 751 -233 757 -199
rect 791 -233 797 -199
rect 751 -271 797 -233
rect 751 -305 757 -271
rect 791 -305 797 -271
rect 751 -343 797 -305
rect 751 -377 757 -343
rect 791 -377 797 -343
rect 751 -415 797 -377
rect 751 -449 757 -415
rect 791 -449 797 -415
rect 751 -487 797 -449
rect 751 -521 757 -487
rect 791 -521 797 -487
rect 751 -559 797 -521
rect 751 -593 757 -559
rect 791 -593 797 -559
rect 751 -631 797 -593
rect 751 -665 757 -631
rect 791 -665 797 -631
rect 751 -703 797 -665
rect 751 -737 757 -703
rect 791 -737 797 -703
rect 751 -775 797 -737
rect 751 -809 757 -775
rect 791 -809 797 -775
rect 751 -847 797 -809
rect 751 -881 757 -847
rect 791 -881 797 -847
rect 751 -919 797 -881
rect 751 -953 757 -919
rect 791 -953 797 -919
rect 751 -991 797 -953
rect 751 -1025 757 -991
rect 791 -1025 797 -991
rect 751 -1063 797 -1025
rect 751 -1097 757 -1063
rect 791 -1097 797 -1063
rect 751 -1135 797 -1097
rect 751 -1169 757 -1135
rect 791 -1169 797 -1135
rect 751 -1207 797 -1169
rect 751 -1241 757 -1207
rect 791 -1241 797 -1207
rect 751 -1279 797 -1241
rect 751 -1313 757 -1279
rect 791 -1313 797 -1279
rect 751 -1351 797 -1313
rect 751 -1385 757 -1351
rect 791 -1385 797 -1351
rect 751 -1423 797 -1385
rect 751 -1457 757 -1423
rect 791 -1457 797 -1423
rect 751 -1495 797 -1457
rect 751 -1529 757 -1495
rect 791 -1529 797 -1495
rect 751 -1567 797 -1529
rect 751 -1601 757 -1567
rect 791 -1601 797 -1567
rect 751 -1639 797 -1601
rect 751 -1673 757 -1639
rect 791 -1673 797 -1639
rect 751 -1711 797 -1673
rect 751 -1745 757 -1711
rect 791 -1745 797 -1711
rect 751 -1783 797 -1745
rect 751 -1817 757 -1783
rect 791 -1817 797 -1783
rect 751 -1855 797 -1817
rect 751 -1889 757 -1855
rect 791 -1889 797 -1855
rect 751 -1927 797 -1889
rect 751 -1961 757 -1927
rect 791 -1961 797 -1927
rect 751 -1999 797 -1961
rect 751 -2033 757 -1999
rect 791 -2033 797 -1999
rect 751 -2071 797 -2033
rect 751 -2105 757 -2071
rect 791 -2105 797 -2071
rect 751 -2143 797 -2105
rect 751 -2177 757 -2143
rect 791 -2177 797 -2143
rect 751 -2215 797 -2177
rect 751 -2249 757 -2215
rect 791 -2249 797 -2215
rect 751 -2287 797 -2249
rect 751 -2321 757 -2287
rect 791 -2321 797 -2287
rect 751 -2359 797 -2321
rect 751 -2393 757 -2359
rect 791 -2393 797 -2359
rect 751 -2431 797 -2393
rect 751 -2465 757 -2431
rect 791 -2465 797 -2431
rect 751 -2500 797 -2465
rect 1009 2465 1055 2500
rect 1009 2431 1015 2465
rect 1049 2431 1055 2465
rect 1009 2393 1055 2431
rect 1009 2359 1015 2393
rect 1049 2359 1055 2393
rect 1009 2321 1055 2359
rect 1009 2287 1015 2321
rect 1049 2287 1055 2321
rect 1009 2249 1055 2287
rect 1009 2215 1015 2249
rect 1049 2215 1055 2249
rect 1009 2177 1055 2215
rect 1009 2143 1015 2177
rect 1049 2143 1055 2177
rect 1009 2105 1055 2143
rect 1009 2071 1015 2105
rect 1049 2071 1055 2105
rect 1009 2033 1055 2071
rect 1009 1999 1015 2033
rect 1049 1999 1055 2033
rect 1009 1961 1055 1999
rect 1009 1927 1015 1961
rect 1049 1927 1055 1961
rect 1009 1889 1055 1927
rect 1009 1855 1015 1889
rect 1049 1855 1055 1889
rect 1009 1817 1055 1855
rect 1009 1783 1015 1817
rect 1049 1783 1055 1817
rect 1009 1745 1055 1783
rect 1009 1711 1015 1745
rect 1049 1711 1055 1745
rect 1009 1673 1055 1711
rect 1009 1639 1015 1673
rect 1049 1639 1055 1673
rect 1009 1601 1055 1639
rect 1009 1567 1015 1601
rect 1049 1567 1055 1601
rect 1009 1529 1055 1567
rect 1009 1495 1015 1529
rect 1049 1495 1055 1529
rect 1009 1457 1055 1495
rect 1009 1423 1015 1457
rect 1049 1423 1055 1457
rect 1009 1385 1055 1423
rect 1009 1351 1015 1385
rect 1049 1351 1055 1385
rect 1009 1313 1055 1351
rect 1009 1279 1015 1313
rect 1049 1279 1055 1313
rect 1009 1241 1055 1279
rect 1009 1207 1015 1241
rect 1049 1207 1055 1241
rect 1009 1169 1055 1207
rect 1009 1135 1015 1169
rect 1049 1135 1055 1169
rect 1009 1097 1055 1135
rect 1009 1063 1015 1097
rect 1049 1063 1055 1097
rect 1009 1025 1055 1063
rect 1009 991 1015 1025
rect 1049 991 1055 1025
rect 1009 953 1055 991
rect 1009 919 1015 953
rect 1049 919 1055 953
rect 1009 881 1055 919
rect 1009 847 1015 881
rect 1049 847 1055 881
rect 1009 809 1055 847
rect 1009 775 1015 809
rect 1049 775 1055 809
rect 1009 737 1055 775
rect 1009 703 1015 737
rect 1049 703 1055 737
rect 1009 665 1055 703
rect 1009 631 1015 665
rect 1049 631 1055 665
rect 1009 593 1055 631
rect 1009 559 1015 593
rect 1049 559 1055 593
rect 1009 521 1055 559
rect 1009 487 1015 521
rect 1049 487 1055 521
rect 1009 449 1055 487
rect 1009 415 1015 449
rect 1049 415 1055 449
rect 1009 377 1055 415
rect 1009 343 1015 377
rect 1049 343 1055 377
rect 1009 305 1055 343
rect 1009 271 1015 305
rect 1049 271 1055 305
rect 1009 233 1055 271
rect 1009 199 1015 233
rect 1049 199 1055 233
rect 1009 161 1055 199
rect 1009 127 1015 161
rect 1049 127 1055 161
rect 1009 89 1055 127
rect 1009 55 1015 89
rect 1049 55 1055 89
rect 1009 17 1055 55
rect 1009 -17 1015 17
rect 1049 -17 1055 17
rect 1009 -55 1055 -17
rect 1009 -89 1015 -55
rect 1049 -89 1055 -55
rect 1009 -127 1055 -89
rect 1009 -161 1015 -127
rect 1049 -161 1055 -127
rect 1009 -199 1055 -161
rect 1009 -233 1015 -199
rect 1049 -233 1055 -199
rect 1009 -271 1055 -233
rect 1009 -305 1015 -271
rect 1049 -305 1055 -271
rect 1009 -343 1055 -305
rect 1009 -377 1015 -343
rect 1049 -377 1055 -343
rect 1009 -415 1055 -377
rect 1009 -449 1015 -415
rect 1049 -449 1055 -415
rect 1009 -487 1055 -449
rect 1009 -521 1015 -487
rect 1049 -521 1055 -487
rect 1009 -559 1055 -521
rect 1009 -593 1015 -559
rect 1049 -593 1055 -559
rect 1009 -631 1055 -593
rect 1009 -665 1015 -631
rect 1049 -665 1055 -631
rect 1009 -703 1055 -665
rect 1009 -737 1015 -703
rect 1049 -737 1055 -703
rect 1009 -775 1055 -737
rect 1009 -809 1015 -775
rect 1049 -809 1055 -775
rect 1009 -847 1055 -809
rect 1009 -881 1015 -847
rect 1049 -881 1055 -847
rect 1009 -919 1055 -881
rect 1009 -953 1015 -919
rect 1049 -953 1055 -919
rect 1009 -991 1055 -953
rect 1009 -1025 1015 -991
rect 1049 -1025 1055 -991
rect 1009 -1063 1055 -1025
rect 1009 -1097 1015 -1063
rect 1049 -1097 1055 -1063
rect 1009 -1135 1055 -1097
rect 1009 -1169 1015 -1135
rect 1049 -1169 1055 -1135
rect 1009 -1207 1055 -1169
rect 1009 -1241 1015 -1207
rect 1049 -1241 1055 -1207
rect 1009 -1279 1055 -1241
rect 1009 -1313 1015 -1279
rect 1049 -1313 1055 -1279
rect 1009 -1351 1055 -1313
rect 1009 -1385 1015 -1351
rect 1049 -1385 1055 -1351
rect 1009 -1423 1055 -1385
rect 1009 -1457 1015 -1423
rect 1049 -1457 1055 -1423
rect 1009 -1495 1055 -1457
rect 1009 -1529 1015 -1495
rect 1049 -1529 1055 -1495
rect 1009 -1567 1055 -1529
rect 1009 -1601 1015 -1567
rect 1049 -1601 1055 -1567
rect 1009 -1639 1055 -1601
rect 1009 -1673 1015 -1639
rect 1049 -1673 1055 -1639
rect 1009 -1711 1055 -1673
rect 1009 -1745 1015 -1711
rect 1049 -1745 1055 -1711
rect 1009 -1783 1055 -1745
rect 1009 -1817 1015 -1783
rect 1049 -1817 1055 -1783
rect 1009 -1855 1055 -1817
rect 1009 -1889 1015 -1855
rect 1049 -1889 1055 -1855
rect 1009 -1927 1055 -1889
rect 1009 -1961 1015 -1927
rect 1049 -1961 1055 -1927
rect 1009 -1999 1055 -1961
rect 1009 -2033 1015 -1999
rect 1049 -2033 1055 -1999
rect 1009 -2071 1055 -2033
rect 1009 -2105 1015 -2071
rect 1049 -2105 1055 -2071
rect 1009 -2143 1055 -2105
rect 1009 -2177 1015 -2143
rect 1049 -2177 1055 -2143
rect 1009 -2215 1055 -2177
rect 1009 -2249 1015 -2215
rect 1049 -2249 1055 -2215
rect 1009 -2287 1055 -2249
rect 1009 -2321 1015 -2287
rect 1049 -2321 1055 -2287
rect 1009 -2359 1055 -2321
rect 1009 -2393 1015 -2359
rect 1049 -2393 1055 -2359
rect 1009 -2431 1055 -2393
rect 1009 -2465 1015 -2431
rect 1049 -2465 1055 -2431
rect 1009 -2500 1055 -2465
rect 1267 2465 1313 2500
rect 1267 2431 1273 2465
rect 1307 2431 1313 2465
rect 1267 2393 1313 2431
rect 1267 2359 1273 2393
rect 1307 2359 1313 2393
rect 1267 2321 1313 2359
rect 1267 2287 1273 2321
rect 1307 2287 1313 2321
rect 1267 2249 1313 2287
rect 1267 2215 1273 2249
rect 1307 2215 1313 2249
rect 1267 2177 1313 2215
rect 1267 2143 1273 2177
rect 1307 2143 1313 2177
rect 1267 2105 1313 2143
rect 1267 2071 1273 2105
rect 1307 2071 1313 2105
rect 1267 2033 1313 2071
rect 1267 1999 1273 2033
rect 1307 1999 1313 2033
rect 1267 1961 1313 1999
rect 1267 1927 1273 1961
rect 1307 1927 1313 1961
rect 1267 1889 1313 1927
rect 1267 1855 1273 1889
rect 1307 1855 1313 1889
rect 1267 1817 1313 1855
rect 1267 1783 1273 1817
rect 1307 1783 1313 1817
rect 1267 1745 1313 1783
rect 1267 1711 1273 1745
rect 1307 1711 1313 1745
rect 1267 1673 1313 1711
rect 1267 1639 1273 1673
rect 1307 1639 1313 1673
rect 1267 1601 1313 1639
rect 1267 1567 1273 1601
rect 1307 1567 1313 1601
rect 1267 1529 1313 1567
rect 1267 1495 1273 1529
rect 1307 1495 1313 1529
rect 1267 1457 1313 1495
rect 1267 1423 1273 1457
rect 1307 1423 1313 1457
rect 1267 1385 1313 1423
rect 1267 1351 1273 1385
rect 1307 1351 1313 1385
rect 1267 1313 1313 1351
rect 1267 1279 1273 1313
rect 1307 1279 1313 1313
rect 1267 1241 1313 1279
rect 1267 1207 1273 1241
rect 1307 1207 1313 1241
rect 1267 1169 1313 1207
rect 1267 1135 1273 1169
rect 1307 1135 1313 1169
rect 1267 1097 1313 1135
rect 1267 1063 1273 1097
rect 1307 1063 1313 1097
rect 1267 1025 1313 1063
rect 1267 991 1273 1025
rect 1307 991 1313 1025
rect 1267 953 1313 991
rect 1267 919 1273 953
rect 1307 919 1313 953
rect 1267 881 1313 919
rect 1267 847 1273 881
rect 1307 847 1313 881
rect 1267 809 1313 847
rect 1267 775 1273 809
rect 1307 775 1313 809
rect 1267 737 1313 775
rect 1267 703 1273 737
rect 1307 703 1313 737
rect 1267 665 1313 703
rect 1267 631 1273 665
rect 1307 631 1313 665
rect 1267 593 1313 631
rect 1267 559 1273 593
rect 1307 559 1313 593
rect 1267 521 1313 559
rect 1267 487 1273 521
rect 1307 487 1313 521
rect 1267 449 1313 487
rect 1267 415 1273 449
rect 1307 415 1313 449
rect 1267 377 1313 415
rect 1267 343 1273 377
rect 1307 343 1313 377
rect 1267 305 1313 343
rect 1267 271 1273 305
rect 1307 271 1313 305
rect 1267 233 1313 271
rect 1267 199 1273 233
rect 1307 199 1313 233
rect 1267 161 1313 199
rect 1267 127 1273 161
rect 1307 127 1313 161
rect 1267 89 1313 127
rect 1267 55 1273 89
rect 1307 55 1313 89
rect 1267 17 1313 55
rect 1267 -17 1273 17
rect 1307 -17 1313 17
rect 1267 -55 1313 -17
rect 1267 -89 1273 -55
rect 1307 -89 1313 -55
rect 1267 -127 1313 -89
rect 1267 -161 1273 -127
rect 1307 -161 1313 -127
rect 1267 -199 1313 -161
rect 1267 -233 1273 -199
rect 1307 -233 1313 -199
rect 1267 -271 1313 -233
rect 1267 -305 1273 -271
rect 1307 -305 1313 -271
rect 1267 -343 1313 -305
rect 1267 -377 1273 -343
rect 1307 -377 1313 -343
rect 1267 -415 1313 -377
rect 1267 -449 1273 -415
rect 1307 -449 1313 -415
rect 1267 -487 1313 -449
rect 1267 -521 1273 -487
rect 1307 -521 1313 -487
rect 1267 -559 1313 -521
rect 1267 -593 1273 -559
rect 1307 -593 1313 -559
rect 1267 -631 1313 -593
rect 1267 -665 1273 -631
rect 1307 -665 1313 -631
rect 1267 -703 1313 -665
rect 1267 -737 1273 -703
rect 1307 -737 1313 -703
rect 1267 -775 1313 -737
rect 1267 -809 1273 -775
rect 1307 -809 1313 -775
rect 1267 -847 1313 -809
rect 1267 -881 1273 -847
rect 1307 -881 1313 -847
rect 1267 -919 1313 -881
rect 1267 -953 1273 -919
rect 1307 -953 1313 -919
rect 1267 -991 1313 -953
rect 1267 -1025 1273 -991
rect 1307 -1025 1313 -991
rect 1267 -1063 1313 -1025
rect 1267 -1097 1273 -1063
rect 1307 -1097 1313 -1063
rect 1267 -1135 1313 -1097
rect 1267 -1169 1273 -1135
rect 1307 -1169 1313 -1135
rect 1267 -1207 1313 -1169
rect 1267 -1241 1273 -1207
rect 1307 -1241 1313 -1207
rect 1267 -1279 1313 -1241
rect 1267 -1313 1273 -1279
rect 1307 -1313 1313 -1279
rect 1267 -1351 1313 -1313
rect 1267 -1385 1273 -1351
rect 1307 -1385 1313 -1351
rect 1267 -1423 1313 -1385
rect 1267 -1457 1273 -1423
rect 1307 -1457 1313 -1423
rect 1267 -1495 1313 -1457
rect 1267 -1529 1273 -1495
rect 1307 -1529 1313 -1495
rect 1267 -1567 1313 -1529
rect 1267 -1601 1273 -1567
rect 1307 -1601 1313 -1567
rect 1267 -1639 1313 -1601
rect 1267 -1673 1273 -1639
rect 1307 -1673 1313 -1639
rect 1267 -1711 1313 -1673
rect 1267 -1745 1273 -1711
rect 1307 -1745 1313 -1711
rect 1267 -1783 1313 -1745
rect 1267 -1817 1273 -1783
rect 1307 -1817 1313 -1783
rect 1267 -1855 1313 -1817
rect 1267 -1889 1273 -1855
rect 1307 -1889 1313 -1855
rect 1267 -1927 1313 -1889
rect 1267 -1961 1273 -1927
rect 1307 -1961 1313 -1927
rect 1267 -1999 1313 -1961
rect 1267 -2033 1273 -1999
rect 1307 -2033 1313 -1999
rect 1267 -2071 1313 -2033
rect 1267 -2105 1273 -2071
rect 1307 -2105 1313 -2071
rect 1267 -2143 1313 -2105
rect 1267 -2177 1273 -2143
rect 1307 -2177 1313 -2143
rect 1267 -2215 1313 -2177
rect 1267 -2249 1273 -2215
rect 1307 -2249 1313 -2215
rect 1267 -2287 1313 -2249
rect 1267 -2321 1273 -2287
rect 1307 -2321 1313 -2287
rect 1267 -2359 1313 -2321
rect 1267 -2393 1273 -2359
rect 1307 -2393 1313 -2359
rect 1267 -2431 1313 -2393
rect 1267 -2465 1273 -2431
rect 1307 -2465 1313 -2431
rect 1267 -2500 1313 -2465
rect -1257 -2538 -1065 -2532
rect -1257 -2572 -1214 -2538
rect -1180 -2572 -1142 -2538
rect -1108 -2572 -1065 -2538
rect -1257 -2578 -1065 -2572
rect -999 -2538 -807 -2532
rect -999 -2572 -956 -2538
rect -922 -2572 -884 -2538
rect -850 -2572 -807 -2538
rect -999 -2578 -807 -2572
rect -741 -2538 -549 -2532
rect -741 -2572 -698 -2538
rect -664 -2572 -626 -2538
rect -592 -2572 -549 -2538
rect -741 -2578 -549 -2572
rect -483 -2538 -291 -2532
rect -483 -2572 -440 -2538
rect -406 -2572 -368 -2538
rect -334 -2572 -291 -2538
rect -483 -2578 -291 -2572
rect -225 -2538 -33 -2532
rect -225 -2572 -182 -2538
rect -148 -2572 -110 -2538
rect -76 -2572 -33 -2538
rect -225 -2578 -33 -2572
rect 33 -2538 225 -2532
rect 33 -2572 76 -2538
rect 110 -2572 148 -2538
rect 182 -2572 225 -2538
rect 33 -2578 225 -2572
rect 291 -2538 483 -2532
rect 291 -2572 334 -2538
rect 368 -2572 406 -2538
rect 440 -2572 483 -2538
rect 291 -2578 483 -2572
rect 549 -2538 741 -2532
rect 549 -2572 592 -2538
rect 626 -2572 664 -2538
rect 698 -2572 741 -2538
rect 549 -2578 741 -2572
rect 807 -2538 999 -2532
rect 807 -2572 850 -2538
rect 884 -2572 922 -2538
rect 956 -2572 999 -2538
rect 807 -2578 999 -2572
rect 1065 -2538 1257 -2532
rect 1065 -2572 1108 -2538
rect 1142 -2572 1180 -2538
rect 1214 -2572 1257 -2538
rect 1065 -2578 1257 -2572
<< properties >>
string FIXED_BBOX -1404 -2657 1404 2657
<< end >>
