* NGSPICE file created from inv_sky130_a_v4.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_L9KS9E a_n73_n81# a_n175_n193# a_n33_41# a_15_n81#
X0 a_15_n81# a_n33_41# a_n73_n81# a_n175_n193# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
**devattr s=5800,316 d=5800,316
C0 a_n33_41# a_n73_n81# 0.014409f
C1 a_n73_n81# a_15_n81# 0.083854f
C2 a_n33_41# a_15_n81# 0.014409f
C3 a_15_n81# a_n175_n193# 0.088419f
C4 a_n73_n81# a_n175_n193# 0.088419f
C5 a_n33_41# a_n175_n193# 0.227f
.ends

.subckt sky130_fd_pr__nfet_01v8_4MHCRP a_2029_n2500# a_n4247_n2674# a_n2029_n2588#
+ a_29_n2588# a_4087_n2500# a_n29_n2500# a_n2087_n2500# a_2087_n2588# a_n4087_n2588#
+ a_n4145_n2500#
X0 a_4087_n2500# a_2087_n2588# a_2029_n2500# a_n4247_n2674# sky130_fd_pr__nfet_01v8 ad=7.25 pd=50.58 as=3.625 ps=25.29 w=25 l=10
**devattr s=145000,5058 d=290000,10116
X1 a_n29_n2500# a_n2029_n2588# a_n2087_n2500# a_n4247_n2674# sky130_fd_pr__nfet_01v8 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=10
**devattr s=145000,5058 d=145000,5058
X2 a_2029_n2500# a_29_n2588# a_n29_n2500# a_n4247_n2674# sky130_fd_pr__nfet_01v8 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=10
**devattr s=145000,5058 d=145000,5058
X3 a_n2087_n2500# a_n4087_n2588# a_n4145_n2500# a_n4247_n2674# sky130_fd_pr__nfet_01v8 ad=3.625 pd=25.29 as=7.25 ps=50.58 w=25 l=10
**devattr s=290000,10116 d=145000,5058
C0 a_n4087_n2588# a_n2029_n2588# 0.104496f
C1 a_2087_n2588# a_4087_n2500# 1.36078f
C2 a_2087_n2588# a_2029_n2500# 1.36078f
C3 a_29_n2588# a_2029_n2500# 1.36078f
C4 a_29_n2588# a_n29_n2500# 1.36078f
C5 a_29_n2588# a_2087_n2588# 0.104496f
C6 a_n2029_n2588# a_n29_n2500# 1.36078f
C7 a_n2029_n2588# a_n2087_n2500# 1.36078f
C8 a_n4087_n2588# a_n2087_n2500# 1.36078f
C9 a_n4087_n2588# a_n4145_n2500# 1.36078f
C10 a_n2029_n2588# a_29_n2588# 0.104496f
C11 a_4087_n2500# a_n4247_n2674# 3.45927f
C12 a_2029_n2500# a_n4247_n2674# 1.88354f
C13 a_n29_n2500# a_n4247_n2674# 1.88016f
C14 a_n2087_n2500# a_n4247_n2674# 1.88354f
C15 a_n4145_n2500# a_n4247_n2674# 3.45927f
C16 a_2087_n2588# a_n4247_n2674# 6.22045f
C17 a_29_n2588# a_n4247_n2674# 6.14529f
C18 a_n2029_n2588# a_n4247_n2674# 6.14529f
C19 a_n4087_n2588# a_n4247_n2674# 6.22045f
.ends

.subckt sky130_fd_pr__nfet_01v8_FPTJ7W a_n1261_n2588# a_n1319_n2500# a_287_n2588#
+ a_487_n2500# a_n287_n2500# a_545_n2588# a_29_n2588# a_n487_n2588# a_745_n2500# a_n545_n2500#
+ a_1003_n2500# a_n29_n2500# a_803_n2588# a_n745_n2588# a_n1003_n2588# a_229_n2500#
+ a_n803_n2500# a_n1421_n2674# a_n229_n2588# a_1261_n2500# a_n1061_n2500# a_1061_n2588#
X0 a_487_n2500# a_287_n2588# a_229_n2500# a_n1421_n2674# sky130_fd_pr__nfet_01v8 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
**devattr s=145000,5058 d=145000,5058
X1 a_n287_n2500# a_n487_n2588# a_n545_n2500# a_n1421_n2674# sky130_fd_pr__nfet_01v8 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
**devattr s=145000,5058 d=145000,5058
X2 a_n29_n2500# a_n229_n2588# a_n287_n2500# a_n1421_n2674# sky130_fd_pr__nfet_01v8 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
**devattr s=145000,5058 d=145000,5058
X3 a_745_n2500# a_545_n2588# a_487_n2500# a_n1421_n2674# sky130_fd_pr__nfet_01v8 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
**devattr s=145000,5058 d=145000,5058
X4 a_1261_n2500# a_1061_n2588# a_1003_n2500# a_n1421_n2674# sky130_fd_pr__nfet_01v8 ad=7.25 pd=50.58 as=3.625 ps=25.29 w=25 l=1
**devattr s=145000,5058 d=290000,10116
X5 a_n545_n2500# a_n745_n2588# a_n803_n2500# a_n1421_n2674# sky130_fd_pr__nfet_01v8 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
**devattr s=145000,5058 d=145000,5058
X6 a_229_n2500# a_29_n2588# a_n29_n2500# a_n1421_n2674# sky130_fd_pr__nfet_01v8 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
**devattr s=145000,5058 d=145000,5058
X7 a_1003_n2500# a_803_n2588# a_745_n2500# a_n1421_n2674# sky130_fd_pr__nfet_01v8 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
**devattr s=145000,5058 d=145000,5058
X8 a_n1061_n2500# a_n1261_n2588# a_n1319_n2500# a_n1421_n2674# sky130_fd_pr__nfet_01v8 ad=3.625 pd=25.29 as=7.25 ps=50.58 w=25 l=1
**devattr s=290000,10116 d=145000,5058
X9 a_n803_n2500# a_n1003_n2588# a_n1061_n2500# a_n1421_n2674# sky130_fd_pr__nfet_01v8 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
**devattr s=145000,5058 d=145000,5058
C0 a_n29_n2500# a_229_n2500# 1.3782f
C1 a_1061_n2588# a_1261_n2500# 0.759836f
C2 a_n287_n2500# a_n29_n2500# 1.3782f
C3 a_1061_n2588# a_1003_n2500# 0.759836f
C4 a_803_n2588# a_1003_n2500# 0.759836f
C5 a_n545_n2500# a_n287_n2500# 1.3782f
C6 a_803_n2588# a_745_n2500# 0.759836f
C7 a_n803_n2500# a_n545_n2500# 1.3782f
C8 a_545_n2588# a_745_n2500# 0.759836f
C9 a_545_n2588# a_487_n2500# 0.759836f
C10 a_n1061_n2500# a_n803_n2500# 1.3782f
C11 a_287_n2588# a_487_n2500# 0.759836f
C12 a_287_n2588# a_229_n2500# 0.759836f
C13 a_n1319_n2500# a_n1061_n2500# 1.3782f
C14 a_29_n2588# a_229_n2500# 0.759836f
C15 a_29_n2588# a_n29_n2500# 0.759836f
C16 a_n229_n2588# a_n29_n2500# 0.759836f
C17 a_n229_n2588# a_n287_n2500# 0.759836f
C18 a_n1261_n2588# a_n1003_n2588# 0.104496f
C19 a_803_n2588# a_1061_n2588# 0.104496f
C20 a_n487_n2588# a_n287_n2500# 0.759836f
C21 a_n487_n2588# a_n545_n2500# 0.759836f
C22 a_545_n2588# a_803_n2588# 0.104496f
C23 a_n745_n2588# a_n545_n2500# 0.759836f
C24 a_n745_n2588# a_n803_n2500# 0.759836f
C25 a_287_n2588# a_545_n2588# 0.104496f
C26 a_29_n2588# a_287_n2588# 0.104496f
C27 a_n229_n2588# a_29_n2588# 0.104496f
C28 a_n487_n2588# a_n229_n2588# 0.104496f
C29 a_n745_n2588# a_n487_n2588# 0.104496f
C30 a_n1003_n2588# a_n803_n2500# 0.759836f
C31 a_n1003_n2588# a_n1061_n2500# 0.759836f
C32 a_n1261_n2588# a_n1061_n2500# 0.759836f
C33 a_n1261_n2588# a_n1319_n2500# 0.759836f
C34 a_n1003_n2588# a_n745_n2588# 0.104496f
C35 a_1003_n2500# a_1261_n2500# 1.3782f
C36 a_745_n2500# a_1003_n2500# 1.3782f
C37 a_487_n2500# a_745_n2500# 1.3782f
C38 a_229_n2500# a_487_n2500# 1.3782f
C39 a_1261_n2500# a_n1421_n2674# 2.812f
C40 a_1003_n2500# a_n1421_n2674# 0.589001f
C41 a_745_n2500# a_n1421_n2674# 0.5881f
C42 a_487_n2500# a_n1421_n2674# 0.587649f
C43 a_229_n2500# a_n1421_n2674# 0.589001f
C44 a_n29_n2500# a_n1421_n2674# 0.592373f
C45 a_n287_n2500# a_n1421_n2674# 0.589001f
C46 a_n545_n2500# a_n1421_n2674# 0.587649f
C47 a_n803_n2500# a_n1421_n2674# 0.5881f
C48 a_n1061_n2500# a_n1421_n2674# 0.589001f
C49 a_n1319_n2500# a_n1421_n2674# 2.812f
C50 a_1061_n2588# a_n1421_n2674# 0.688382f
C51 a_803_n2588# a_n1421_n2674# 0.619772f
C52 a_545_n2588# a_n1421_n2674# 0.618982f
C53 a_287_n2588# a_n1421_n2674# 0.618685f
C54 a_29_n2588# a_n1421_n2674# 0.618449f
C55 a_n229_n2588# a_n1421_n2674# 0.618449f
C56 a_n487_n2588# a_n1421_n2674# 0.618685f
C57 a_n745_n2588# a_n1421_n2674# 0.618982f
C58 a_n1003_n2588# a_n1421_n2674# 0.619772f
C59 a_n1261_n2588# a_n1421_n2674# 0.688382f
.ends

.subckt sky130_fd_pr__pfet_01v8_ND7MJ4 a_79_n2500# a_295_n2500# a_n411_n2597# a_187_n2500#
+ a_21_n2597# a_n461_n2500# a_237_n2597# a_n353_n2500# a_345_2531# a_129_2531# a_n245_n2500#
+ a_n29_n2500# a_n137_n2500# a_n195_n2597# w_n599_n2719# a_403_n2500# a_n87_2531#
+ a_n303_2531# VSUBS
X0 a_n353_n2500# a_n411_n2597# a_n461_n2500# w_n599_n2719# sky130_fd_pr__pfet_01v8 ad=3.625 pd=25.29 as=7.25 ps=50.58 w=25 l=0.25
**devattr s=290000,10116 d=145000,5058
X1 a_187_n2500# a_129_2531# a_79_n2500# w_n599_n2719# sky130_fd_pr__pfet_01v8 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=0.25
**devattr s=145000,5058 d=145000,5058
X2 a_n137_n2500# a_n195_n2597# a_n245_n2500# w_n599_n2719# sky130_fd_pr__pfet_01v8 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=0.25
**devattr s=145000,5058 d=145000,5058
X3 a_n29_n2500# a_n87_2531# a_n137_n2500# w_n599_n2719# sky130_fd_pr__pfet_01v8 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=0.25
**devattr s=145000,5058 d=145000,5058
X4 a_79_n2500# a_21_n2597# a_n29_n2500# w_n599_n2719# sky130_fd_pr__pfet_01v8 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=0.25
**devattr s=145000,5058 d=145000,5058
X5 a_295_n2500# a_237_n2597# a_187_n2500# w_n599_n2719# sky130_fd_pr__pfet_01v8 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=0.25
**devattr s=145000,5058 d=145000,5058
X6 a_n245_n2500# a_n303_2531# a_n353_n2500# w_n599_n2719# sky130_fd_pr__pfet_01v8 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=0.25
**devattr s=145000,5058 d=145000,5058
X7 a_403_n2500# a_345_2531# a_295_n2500# w_n599_n2719# sky130_fd_pr__pfet_01v8 ad=7.25 pd=50.58 as=3.625 ps=25.29 w=25 l=0.25
**devattr s=145000,5058 d=290000,10116
C0 a_187_n2500# a_295_n2500# 3.27775f
C1 a_79_n2500# a_187_n2500# 3.27775f
C2 a_n29_n2500# a_79_n2500# 3.27775f
C3 a_n137_n2500# a_n29_n2500# 3.27775f
C4 a_237_n2597# a_295_n2500# 0.259865f
C5 a_n245_n2500# a_n137_n2500# 3.27775f
C6 a_237_n2597# a_187_n2500# 0.259865f
C7 a_n353_n2500# a_n245_n2500# 3.27775f
C8 a_21_n2597# a_79_n2500# 0.259865f
C9 a_345_2531# a_403_n2500# 0.259865f
C10 a_21_n2597# a_n29_n2500# 0.259865f
C11 a_345_2531# a_295_n2500# 0.259865f
C12 a_n461_n2500# a_n353_n2500# 3.27775f
C13 a_n195_n2597# a_n137_n2500# 0.259865f
C14 a_129_2531# a_187_n2500# 0.259865f
C15 w_n599_n2719# a_n303_2531# 0.127054f
C16 a_n195_n2597# a_n245_n2500# 0.259865f
C17 a_129_2531# a_79_n2500# 0.259865f
C18 a_21_n2597# a_237_n2597# 0.022307f
C19 a_n411_n2597# a_n353_n2500# 0.259865f
C20 a_n87_2531# a_n29_n2500# 0.259865f
C21 a_n411_n2597# a_n461_n2500# 0.259865f
C22 a_n87_2531# a_n137_n2500# 0.259865f
C23 a_n195_n2597# a_21_n2597# 0.022307f
C24 a_345_2531# a_237_n2597# 0.014345f
C25 a_n411_n2597# a_n195_n2597# 0.022307f
C26 a_129_2531# a_237_n2597# 0.014345f
C27 a_129_2531# a_21_n2597# 0.014345f
C28 a_n87_2531# a_21_n2597# 0.014345f
C29 a_n87_2531# a_n195_n2597# 0.014345f
C30 a_129_2531# a_345_2531# 0.022307f
C31 a_n87_2531# a_129_2531# 0.022307f
C32 w_n599_n2719# a_403_n2500# 1.62409f
C33 w_n599_n2719# a_295_n2500# 0.023582f
C34 w_n599_n2719# a_187_n2500# 0.023582f
C35 w_n599_n2719# a_79_n2500# 0.024232f
C36 w_n599_n2719# a_n29_n2500# 0.021322f
C37 w_n599_n2719# a_n137_n2500# 0.024232f
C38 a_n303_2531# a_n245_n2500# 0.259865f
C39 w_n599_n2719# a_n245_n2500# 0.023582f
C40 a_n303_2531# a_n353_n2500# 0.259865f
C41 w_n599_n2719# a_n353_n2500# 0.023582f
C42 w_n599_n2719# a_n461_n2500# 1.62409f
C43 w_n599_n2719# a_237_n2597# 0.127054f
C44 a_n303_2531# a_n195_n2597# 0.014345f
C45 w_n599_n2719# a_21_n2597# 0.116573f
C46 a_n303_2531# a_n411_n2597# 0.014345f
C47 w_n599_n2719# a_n195_n2597# 0.115341f
C48 w_n599_n2719# a_n411_n2597# 0.130912f
C49 w_n599_n2719# a_345_2531# 0.130912f
C50 a_n303_2531# a_n87_2531# 0.022307f
C51 w_n599_n2719# a_129_2531# 0.115341f
C52 w_n599_n2719# a_n87_2531# 0.116573f
C53 a_295_n2500# a_403_n2500# 3.27775f
C54 a_403_n2500# VSUBS 1.01166f
C55 a_295_n2500# VSUBS 0.218985f
C56 a_187_n2500# VSUBS 0.218985f
C57 a_79_n2500# VSUBS 0.218985f
C58 a_n29_n2500# VSUBS 0.218985f
C59 a_n137_n2500# VSUBS 0.218985f
C60 a_n245_n2500# VSUBS 0.218985f
C61 a_n353_n2500# VSUBS 0.218985f
C62 a_n461_n2500# VSUBS 1.01166f
C63 a_237_n2597# VSUBS 0.068093f
C64 a_21_n2597# VSUBS 0.058829f
C65 a_n195_n2597# VSUBS 0.058829f
C66 a_n411_n2597# VSUBS 0.07532f
C67 a_345_2531# VSUBS 0.07532f
C68 a_129_2531# VSUBS 0.058829f
C69 a_n87_2531# VSUBS 0.058829f
C70 a_n303_2531# VSUBS 0.068093f
C71 w_n599_n2719# VSUBS 22.3107f
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_5UY5E6 m3_n2786_n2640# c1_n2746_n2600# VSUBS
X0 c1_n2746_n2600# m3_n2786_n2640# sky130_fd_pr__cap_mim_m3_1 l=26 w=26
C0 m3_n2786_n2640# c1_n2746_n2600# 59.715103f
C1 c1_n2746_n2600# VSUBS 2.69897f
C2 m3_n2786_n2640# VSUBS 14.5533f
.ends

.subckt inv_sky130_a_v4 VG1 VCC VG2 out in VSS
XXM1 m1_8420_9480# VSS VG1 m1_6370_6630# sky130_fd_pr__nfet_01v8_L9KS9E
XXM3 VSS VSS out out VSS VSS VSS out out VSS sky130_fd_pr__nfet_01v8_4MHCRP
XXM4 m1_6370_6630# m1_8420_9480# m1_6370_6630# VSS m1_8420_9480# m1_6370_6630# m1_6370_6630#
+ m1_6370_6630# m1_8420_9480# VSS VSS VSS m1_6370_6630# m1_6370_6630# m1_6370_6630#
+ m1_8420_9480# m1_8420_9480# VSS m1_6370_6630# m1_8420_9480# VSS m1_6370_6630# sky130_fd_pr__nfet_01v8_FPTJ7W
XXM5 m1_8420_9480# m1_8420_9480# m1_6370_6630# VCC m1_6370_6630# VCC m1_6370_6630#
+ m1_8420_9480# m1_6370_6630# m1_6370_6630# VCC VCC m1_8420_9480# m1_6370_6630# VCC
+ VCC m1_6370_6630# m1_6370_6630# VSS sky130_fd_pr__pfet_01v8_ND7MJ4
XXC1 m1_6370_6630# in VSS sky130_fd_pr__cap_mim_m3_1_5UY5E6
Xsky130_fd_pr__nfet_01v8_L9KS9E_0 m1_8420_9480# VSS VG2 out sky130_fd_pr__nfet_01v8_L9KS9E
C0 VG1 VG2 9.11e-19
C1 VG1 in -9.16e-35
C2 VCC VG2 0.019075f
C3 out m1_6370_6630# 12.586376f
C4 m1_8420_9480# VG2 0.130126f
C5 m1_8420_9480# in -2.73e-32
C6 VG1 VCC 0.018291f
C7 m1_6370_6630# VG2 0.220862f
C8 m1_6370_6630# in 0.188818f
C9 VG1 m1_8420_9480# 0.106703f
C10 m1_8420_9480# VCC 1.632583f
C11 out VG2 0.052763f
C12 out in 1.179613f
C13 VG1 m1_6370_6630# 0.223186f
C14 m1_6370_6630# VCC 5.088756f
C15 VG1 out 0.001196f
C16 m1_6370_6630# m1_8420_9480# 10.49333f
C17 in VG2 9.16e-35
C18 out m1_8420_9480# 0.665724f
C19 VG2 VSS 0.431946f
C20 in VSS 2.908484f
C21 VCC VSS 24.962215f
C22 m1_8420_9480# VSS 12.487506f
C23 m1_6370_6630# VSS 35.560314f
C24 out VSS 37.053707f
C25 VG1 VSS 0.414288f
.ends

