** sch_path: /Users/miguelcorrea/Desktop/MA2_project/Amplifier_Inv/xschem/biasing_test.sch
**.subckt biasing_test
x1 out in VCC VSS not W_N=20 L_N=0.15 W_P=40 L_P=0.15 m=1
VN VSS GND 0
VP VCC GND 1.5
Vin in GND 0.7052
C1 out GND 1p m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt




.control
  op
  print @m.x1.xm1.msky130_fd_pr__nfet_01v8[gm]
  print @m.x1.xm2.msky130_fd_pr__pfet_01v8[gm]
  print @m.x1.xm1.msky130_fd_pr__nfet_01v8[gds]
  print @m.x1.xm2.msky130_fd_pr__pfet_01v8[gds]
  print @m.x1.xm1.msky130_fd_pr__nfet_01v8[cgs]
  print @m.x1.xm2.msky130_fd_pr__pfet_01v8[cgs]
  save all
  write tb_inv_sky130_op.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  sky130_tests/not.sym # of pins=2
** sym_path: /usr/local/share/pdk/sky130A/libs.tech/xschem/sky130_tests/not.sym
** sch_path: /usr/local/share/pdk/sky130A/libs.tech/xschem/sky130_tests/not.sch
.subckt not y a VCCPIN VSSPIN     W_N=1 L_N=0.15 W_P=2 L_P=0.15
*.opin y
*.ipin a
XM1 y a VSSPIN VSSPIN sky130_fd_pr__nfet_01v8 L=L_N W=W_N nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 y a VCCPIN VCCPIN sky130_fd_pr__pfet_01v8 L=L_P W=W_P nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.GLOBAL VSS
.GLOBAL VCC
.end
