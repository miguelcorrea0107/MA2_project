magic
tech sky130A
magscale 1 2
timestamp 1716656893
<< nwell >>
rect 7660 10850 10310 11040
rect 7660 10810 10420 10850
rect 7770 10800 10420 10810
<< pwell >>
rect 9670 9570 9690 9650
rect 6300 9280 11680 9390
rect 6340 9270 11680 9280
rect 7720 6250 10480 6580
<< locali >>
rect 6250 11190 11730 11210
rect 6250 11030 6510 11190
rect 11720 11030 11730 11190
rect 6250 10914 11730 11030
rect 6250 10910 7660 10914
rect 10420 10910 11730 10914
rect 6250 9810 6320 10910
rect 7770 10800 10420 10810
rect 11660 9810 11730 10910
rect 6250 9800 11730 9810
rect 6250 9280 11730 9390
rect 6250 6460 6320 9280
rect 6340 9270 11730 9280
rect 11650 6460 11730 9270
rect 6250 6370 11730 6460
rect 6250 -2100 6320 6370
rect 11650 -2100 11730 6370
rect 6250 -2200 11730 -2100
rect 6250 -2360 6510 -2200
rect 11720 -2360 11730 -2200
rect 6250 -2380 11730 -2360
<< viali >>
rect 6510 11030 11720 11190
rect 6510 -2360 11720 -2200
<< metal1 >>
rect 6250 11190 11730 11210
rect 6250 11030 6510 11190
rect 11720 11030 11730 11190
rect 6250 11010 11730 11030
rect 6370 10710 6380 10780
rect 6450 10710 6460 10780
rect 8880 10770 8890 10832
rect 9210 10770 9220 10832
rect 7554 10664 7564 10726
rect 7884 10664 7894 10726
rect 6370 10500 6380 10570
rect 6450 10500 6460 10570
rect 8880 10552 8890 10614
rect 9210 10552 9220 10614
rect 11520 10610 11530 10670
rect 11590 10610 11600 10670
rect 7552 10440 7562 10502
rect 7882 10440 7892 10502
rect 11520 10400 11530 10460
rect 11590 10400 11600 10460
rect 6370 10280 6380 10350
rect 6450 10280 6460 10350
rect 8880 10336 8890 10398
rect 9210 10336 9220 10398
rect 7552 10222 7562 10284
rect 7882 10222 7892 10284
rect 6370 10060 6380 10130
rect 6450 10060 6460 10130
rect 8880 10120 8890 10182
rect 9210 10120 9220 10182
rect 11520 10180 11530 10240
rect 11590 10180 11600 10240
rect 7552 10012 7562 10074
rect 7882 10012 7892 10074
rect 9560 10020 9570 10074
rect 9690 10020 9700 10074
rect 8880 9910 8890 9972
rect 9210 9910 9220 9972
rect 11520 9960 11530 10020
rect 11590 9960 11600 10020
rect 6370 9780 6380 9880
rect 6460 9780 7170 9880
rect 7370 9870 11520 9880
rect 7370 9800 8420 9870
rect 8510 9800 11520 9870
rect 7370 9780 11520 9800
rect 11590 9780 11600 9880
rect 7980 9590 8280 9650
rect 7980 9520 8380 9590
rect 8410 9580 8420 9650
rect 8510 9580 8520 9650
rect 9560 9645 9570 9650
rect 9265 9595 9570 9645
rect 9265 9530 9315 9595
rect 9560 9580 9570 9595
rect 9670 9580 9680 9650
rect 7980 9450 8280 9520
rect 8420 9480 9315 9530
rect 9570 9400 9580 9520
rect 9670 9400 9680 9520
rect 9710 9460 10110 9660
rect 6370 8950 6380 9130
rect 6440 8950 6450 9130
rect 7548 9124 7558 9196
rect 7880 9124 7890 9196
rect 11510 8950 11520 9130
rect 11580 8950 11590 9130
rect 8670 8878 8680 8940
rect 9000 8878 9010 8940
rect 6370 8690 6380 8870
rect 6440 8690 6450 8870
rect 11510 8690 11520 8870
rect 11580 8690 11590 8870
rect 7552 8616 7562 8678
rect 7882 8616 7892 8678
rect 6370 8430 6380 8610
rect 6440 8430 6450 8610
rect 11510 8430 11520 8610
rect 11580 8430 11590 8610
rect 8664 8360 8674 8422
rect 8994 8360 9004 8422
rect 6370 8170 6380 8350
rect 6440 8170 6450 8350
rect 11510 8170 11520 8350
rect 11580 8170 11590 8350
rect 7550 8098 7560 8160
rect 7880 8098 7890 8160
rect 6370 7910 6380 8090
rect 6440 7910 6450 8090
rect 11510 7910 11520 8090
rect 11580 7910 11590 8090
rect 8668 7846 8678 7908
rect 8998 7846 9008 7908
rect 6370 7660 6380 7840
rect 6440 7660 6450 7840
rect 11510 7660 11520 7840
rect 11580 7660 11590 7840
rect 7552 7584 7562 7646
rect 7882 7584 7892 7646
rect 6370 7400 6380 7580
rect 6440 7400 6450 7580
rect 11510 7400 11520 7580
rect 11580 7400 11590 7580
rect 8670 7326 8680 7388
rect 9000 7326 9010 7388
rect 6370 7140 6380 7320
rect 6440 7140 6450 7320
rect 11510 7140 11520 7320
rect 11580 7140 11590 7320
rect 7556 7068 7566 7130
rect 7886 7068 7896 7130
rect 6370 6880 6380 7060
rect 6440 6880 6450 7060
rect 11510 6880 11520 7060
rect 11580 6880 11590 7060
rect 8668 6814 8678 6876
rect 8998 6814 9008 6876
rect 6370 6630 6380 6810
rect 6440 6630 6450 6810
rect 11510 6630 11520 6810
rect 11580 6630 11590 6810
rect 7554 6552 7564 6614
rect 7884 6552 7894 6614
rect 8672 6222 8682 6284
rect 9002 6222 9012 6284
rect 6370 4230 6380 6210
rect 6440 5960 6450 6210
rect 11510 5960 11520 6220
rect 6440 5940 11520 5960
rect 6440 5640 9580 5940
rect 9660 5640 11520 5940
rect 6440 5620 11520 5640
rect 6440 4230 6450 5620
rect 11510 4230 11520 5620
rect 11580 4230 11590 6220
rect 8674 4158 8684 4220
rect 9004 4158 9014 4220
rect 6370 2170 6380 4150
rect 6440 2170 6450 4150
rect 9670 3684 9680 3884
rect 9880 3684 9890 3884
rect 9680 3484 9880 3684
rect 11510 2170 11520 4160
rect 11580 2170 11590 4160
rect 8668 2102 8678 2164
rect 8998 2102 9008 2164
rect 6370 110 6380 2090
rect 6440 110 6450 2090
rect 11510 110 11520 2100
rect 11580 110 11590 2100
rect 8668 44 8678 106
rect 8998 44 9008 106
rect 6370 -1950 6380 30
rect 6440 -1950 6450 30
rect 11510 -1950 11520 40
rect 11580 -1950 11590 40
rect 8672 -2016 8682 -1954
rect 9002 -2016 9012 -1954
rect 6250 -2198 11730 -2180
rect 6250 -2200 8682 -2198
rect 9008 -2200 11730 -2198
rect 6250 -2360 6510 -2200
rect 11720 -2360 11730 -2200
rect 6250 -2364 8682 -2360
rect 9008 -2364 11730 -2360
rect 6250 -2380 11730 -2364
<< via1 >>
rect 8892 11034 9220 11188
rect 6380 10710 6450 10780
rect 8890 10770 9210 10832
rect 7564 10664 7884 10726
rect 6380 10500 6450 10570
rect 8890 10552 9210 10614
rect 11530 10610 11590 10670
rect 7562 10440 7882 10502
rect 11530 10400 11590 10460
rect 6380 10280 6450 10350
rect 8890 10336 9210 10398
rect 7562 10222 7882 10284
rect 6380 10060 6450 10130
rect 8890 10120 9210 10182
rect 11530 10180 11590 10240
rect 7562 10012 7882 10074
rect 9570 10020 9690 10074
rect 8890 9910 9210 9972
rect 11530 9960 11590 10020
rect 6380 9780 6460 9880
rect 7170 9780 7370 9880
rect 8420 9800 8510 9870
rect 11520 9780 11590 9880
rect 8420 9580 8510 9650
rect 9570 9580 9670 9650
rect 9580 9400 9670 9520
rect 6380 8950 6440 9130
rect 7558 9124 7880 9196
rect 11520 8950 11580 9130
rect 8680 8878 9000 8940
rect 6380 8690 6440 8870
rect 11520 8690 11580 8870
rect 7562 8616 7882 8678
rect 6380 8430 6440 8610
rect 11520 8430 11580 8610
rect 8674 8360 8994 8422
rect 6380 8170 6440 8350
rect 11520 8170 11580 8350
rect 7560 8098 7880 8160
rect 6380 7910 6440 8090
rect 11520 7910 11580 8090
rect 8678 7846 8998 7908
rect 6380 7660 6440 7840
rect 11520 7660 11580 7840
rect 7562 7584 7882 7646
rect 6380 7400 6440 7580
rect 11520 7400 11580 7580
rect 8680 7326 9000 7388
rect 6380 7140 6440 7320
rect 11520 7140 11580 7320
rect 7566 7068 7886 7130
rect 6380 6880 6440 7060
rect 11520 6880 11580 7060
rect 8678 6814 8998 6876
rect 6380 6630 6440 6810
rect 11520 6630 11580 6810
rect 7564 6552 7884 6614
rect 8682 6222 9002 6284
rect 6380 4230 6440 6210
rect 9580 5640 9660 5940
rect 11520 4230 11580 6220
rect 8684 4158 9004 4220
rect 6380 2170 6440 4150
rect 9680 3684 9880 3884
rect 11520 2170 11580 4160
rect 8678 2102 8998 2164
rect 6380 110 6440 2090
rect 11520 110 11580 2100
rect 8678 44 8998 106
rect 6380 -1950 6440 30
rect 11520 -1950 11580 40
rect 8682 -2016 9002 -1954
rect 8682 -2200 9008 -2198
rect 8682 -2360 9008 -2200
rect 8682 -2364 9008 -2360
<< metal2 >>
rect 8892 11190 9220 11198
rect 8890 11188 9220 11190
rect 8890 11034 8892 11188
rect 8890 11024 9220 11034
rect 8890 10832 9210 11024
rect 6370 10780 6470 10790
rect 6370 10710 6380 10780
rect 6450 10710 6470 10780
rect 6370 10570 6470 10710
rect 6370 10500 6380 10570
rect 6450 10500 6470 10570
rect 6370 10350 6470 10500
rect 6370 10280 6380 10350
rect 6450 10280 6470 10350
rect 6370 10130 6470 10280
rect 6370 10060 6380 10130
rect 6450 10060 6470 10130
rect 6370 9880 6470 10060
rect 7562 10736 7882 10746
rect 7562 10726 7884 10736
rect 7562 10664 7564 10726
rect 7562 10654 7884 10664
rect 7562 10502 7882 10654
rect 7562 10284 7882 10440
rect 7562 10074 7882 10222
rect 6370 9780 6380 9880
rect 6460 9780 6470 9880
rect 6370 9130 6470 9780
rect 7170 9880 7370 9890
rect 7170 9770 7370 9780
rect 7180 9560 7360 9770
rect 7180 9470 7360 9480
rect 7562 9206 7882 10012
rect 8890 10614 9210 10770
rect 8890 10398 9210 10552
rect 8890 10182 9210 10336
rect 8890 9972 9210 10120
rect 11510 10670 11600 10780
rect 11510 10610 11530 10670
rect 11590 10610 11600 10670
rect 11510 10460 11600 10610
rect 11510 10400 11530 10460
rect 11590 10400 11600 10460
rect 11510 10240 11600 10400
rect 11510 10180 11530 10240
rect 11590 10180 11600 10240
rect 8890 9898 9210 9910
rect 9570 10074 9690 10094
rect 8420 9870 8510 9880
rect 8420 9650 8510 9800
rect 8420 9570 8510 9580
rect 9570 9650 9690 10020
rect 9670 9580 9690 9650
rect 9570 9570 9690 9580
rect 11510 10020 11600 10180
rect 11510 9960 11530 10020
rect 11590 9960 11600 10020
rect 11510 9880 11600 9960
rect 11510 9780 11520 9880
rect 11590 9780 11600 9880
rect 9580 9520 9670 9530
rect 6370 8950 6380 9130
rect 6440 8950 6470 9130
rect 7558 9196 7882 9206
rect 7880 9124 7882 9196
rect 7558 9114 7882 9124
rect 6370 8870 6470 8950
rect 6370 8690 6380 8870
rect 6440 8690 6470 8870
rect 6370 8610 6470 8690
rect 6370 8430 6380 8610
rect 6440 8430 6470 8610
rect 6370 8350 6470 8430
rect 6370 8170 6380 8350
rect 6440 8170 6470 8350
rect 7562 8678 7882 9114
rect 9570 9400 9580 9520
rect 9670 9400 9680 9520
rect 7562 8170 7882 8616
rect 8680 8940 9000 8978
rect 8680 8432 9000 8878
rect 8674 8422 9000 8432
rect 8994 8360 9000 8422
rect 8674 8350 9000 8360
rect 6370 8090 6470 8170
rect 6370 7910 6380 8090
rect 6440 7910 6470 8090
rect 7560 8160 7882 8170
rect 7880 8098 7882 8160
rect 7560 8088 7882 8098
rect 6370 7840 6470 7910
rect 6370 7660 6380 7840
rect 6440 7660 6470 7840
rect 6370 7580 6470 7660
rect 6370 7400 6380 7580
rect 6440 7400 6470 7580
rect 6370 7320 6470 7400
rect 6370 7140 6380 7320
rect 6440 7140 6470 7320
rect 6370 7060 6470 7140
rect 6370 6880 6380 7060
rect 6440 6880 6470 7060
rect 6370 6810 6470 6880
rect 6370 6630 6380 6810
rect 6440 6630 6470 6810
rect 6370 6610 6470 6630
rect 7562 7646 7882 8088
rect 8680 7918 9000 8350
rect 8678 7908 9000 7918
rect 8998 7846 9000 7908
rect 8678 7836 9000 7846
rect 7562 7140 7882 7584
rect 8680 7388 9000 7836
rect 7562 7130 7886 7140
rect 7562 7068 7566 7130
rect 7562 7058 7886 7068
rect 7562 6624 7882 7058
rect 8680 6886 9000 7326
rect 8678 6876 9000 6886
rect 8998 6814 9000 6876
rect 8678 6804 9000 6814
rect 8680 6656 9000 6804
rect 7562 6614 7884 6624
rect 7562 6552 7564 6614
rect 7562 6546 7884 6552
rect 7564 6542 7884 6546
rect 8680 6476 9002 6656
rect 8682 6284 9002 6476
rect 6370 6210 6450 6230
rect 6370 4230 6380 6210
rect 6440 4230 6450 6210
rect 8682 6066 9002 6222
rect 8680 5840 9002 6066
rect 9570 5940 9680 9400
rect 11510 9130 11600 9780
rect 11510 8950 11520 9130
rect 11580 8950 11600 9130
rect 11510 8870 11600 8950
rect 11510 8690 11520 8870
rect 11580 8690 11600 8870
rect 11510 8610 11600 8690
rect 11510 8430 11520 8610
rect 11580 8430 11600 8610
rect 11510 8350 11600 8430
rect 11510 8170 11520 8350
rect 11580 8170 11600 8350
rect 11510 8090 11600 8170
rect 11510 7910 11520 8090
rect 11580 7910 11600 8090
rect 11510 7840 11600 7910
rect 11510 7660 11520 7840
rect 11580 7660 11600 7840
rect 11510 7580 11600 7660
rect 11510 7400 11520 7580
rect 11580 7400 11600 7580
rect 11510 7320 11600 7400
rect 11510 7140 11520 7320
rect 11580 7140 11600 7320
rect 11510 7060 11600 7140
rect 11510 6880 11520 7060
rect 11580 6880 11600 7060
rect 11510 6810 11600 6880
rect 11510 6630 11520 6810
rect 11580 6630 11600 6810
rect 11510 6610 11600 6630
rect 8680 5620 9000 5840
rect 9570 5640 9580 5940
rect 9660 5640 9680 5940
rect 9570 5620 9680 5640
rect 11500 6220 11590 6240
rect 8680 5250 9002 5620
rect 8682 4904 9002 5250
rect 6370 4150 6450 4230
rect 6370 2170 6380 4150
rect 6440 2170 6450 4150
rect 8680 4804 9002 4904
rect 8680 4230 9000 4804
rect 11500 4230 11520 6220
rect 11580 4230 11590 6220
rect 8680 4220 9004 4230
rect 8680 4158 8684 4220
rect 8680 4148 9004 4158
rect 11500 4160 11590 4230
rect 8680 2174 9000 4148
rect 9680 3884 9880 3894
rect 9680 3674 9880 3684
rect 6370 2090 6450 2170
rect 8678 2164 9000 2174
rect 8998 2102 9000 2164
rect 8678 2092 9000 2102
rect 6370 110 6380 2090
rect 6440 110 6450 2090
rect 8680 116 9000 2092
rect 6370 30 6450 110
rect 8678 106 9000 116
rect 8998 44 9000 106
rect 8678 34 9000 44
rect 6370 -1950 6380 30
rect 6440 -1950 6450 30
rect 8680 -1032 9000 34
rect 11500 2170 11520 4160
rect 11580 2170 11590 4160
rect 11500 2100 11590 2170
rect 11500 110 11520 2100
rect 11580 110 11590 2100
rect 11500 40 11590 110
rect 8680 -1552 9002 -1032
rect 6370 -1970 6450 -1950
rect 8682 -1954 9002 -1552
rect 11500 -1950 11520 40
rect 11580 -1950 11590 40
rect 11500 -1970 11590 -1950
rect 8682 -2188 9002 -2016
rect 8682 -2198 9008 -2188
rect 8682 -2374 9008 -2364
<< via2 >>
rect 7180 9480 7360 9560
rect 9680 3684 9880 3884
<< metal3 >>
rect 9670 3884 9890 3889
rect 9670 3684 9680 3884
rect 9880 3684 9890 3884
rect 9670 3679 9890 3684
<< via3 >>
rect 9680 3684 9880 3884
<< metal4 >>
rect 9680 3885 9880 4138
rect 9679 3884 9881 3885
rect 9679 3684 9680 3884
rect 9880 3684 9881 3884
rect 9679 3683 9881 3684
use sky130_fd_pr__nfet_01v8_L9KS9E  sky130_fd_pr__nfet_01v8_L9KS9E_0
timestamp 1716644424
transform 0 1 9659 -1 0 9551
box -201 -219 201 219
use sky130_fd_pr__cap_mim_m3_1_5UY5E6  XC1
timestamp 1716644424
transform 0 -1 8970 1 0 6786
box -2786 -2640 2786 2640
use sky130_fd_pr__nfet_01v8_L9KS9E  XM1
timestamp 1716644424
transform 0 -1 8429 1 0 9551
box -201 -219 201 219
use sky130_fd_pr__nfet_01v8_4MHCRP  XM3
timestamp 1716644424
transform 0 -1 8980 1 0 2133
box -4273 -2700 4273 2700
use sky130_fd_pr__nfet_01v8_FPTJ7W  XM4
timestamp 1716644424
transform 0 -1 8980 1 0 7877
box -1447 -2700 1447 2700
use sky130_fd_pr__pfet_01v8_ND7MJ4  XM5
timestamp 1716644424
transform 0 1 8989 -1 0 10369
box -599 -2719 599 2719
<< labels >>
flabel metal1 6290 -2380 6490 -2180 0 FreeSans 256 0 0 0 VSS
port 5 nsew
flabel metal1 6290 11010 6490 11210 0 FreeSans 256 0 0 0 VCC
port 1 nsew
flabel metal1 7980 9450 8180 9650 0 FreeSans 256 0 0 0 VG1
port 0 nsew
flabel metal1 9910 9460 10110 9660 0 FreeSans 256 0 0 0 VG2
port 2 nsew
flabel metal1 10310 5730 10510 5930 0 FreeSans 256 0 0 0 out
port 3 nsew
flabel metal1 9680 3484 9880 3684 0 FreeSans 256 0 0 0 in
port 4 nsew
<< end >>
