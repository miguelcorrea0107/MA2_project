** sch_path: /Users/miguelcorrea/Desktop/MA2_project/Amplifier_Inv/xschem/tb_inv_sky130_a.sch
**.subckt tb_inv_sky130_a
VN VSS GND 0
VP VCC GND 1.125
.save i(vp)
Vin in GND 0.44866 ac 1e-3 sin(0.44866 0.001 1000 0 0 0)
.save i(vin)
Rl out GND 1e15 m=1
x1 out in inv_sky130_a
**** begin user architecture code

** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt



.control

  op
  save all
  let gmn = @m.x1.x1.xm1.msky130_fd_pr__nfet_01v8[gm]
  let gmp = @m.x1.x1.xm2.msky130_fd_pr__pfet_01v8[gm]
  let gdsn = @m.x1.x1.xm1.msky130_fd_pr__nfet_01v8[gds]
  let gdsp = @m.x1.x1.xm2.msky130_fd_pr__pfet_01v8[gds]
  let cgsn = @m.x1.x1.xm1.msky130_fd_pr__nfet_01v8[cgs]
  let cgsp = @m.x1.x1.xm2.msky130_fd_pr__pfet_01v8[cgs]
  let vthn = @m.x1.x1.xm1.msky130_fd_pr__nfet_01v8[vth]
  write tb_inv_sky130_a_op.raw gmn gmp gdsn gdsp cgsn cgsp vthn

  ac dec 10000 1 1e5
  save all
  let gain = db(v(out)/v(in))
  let phase = phase(v(out)/v(in))
  write tb_inv_sky130_a_AC.raw gain phase

  noise v(out) Vin dec 1000 300 10k 10
  save all
  write tb_inv_sky130_a_noise.raw

  noise v(out) Vin dec 1000 300 10k
  save all
  setplot noise1
  write tb_inv_sky130_a_noise_spectrum.raw

  tran 0.1u 2m
  save all
  let pw_in = i(Vin)*v(in)
  let pw_vcc = i(Vp)*1,125
  let pw_total = pw_in+pw_vcc
  meas tran avg_pw_total AVG pw_total FROM=0 TO=2m
  meas tran avg_pw_in AVG pw_in FROM=0 TO=2m
  meas tran avg_pw_vcc AVG pw_vcc FROM=0 TO=2m
  write tb_inv_sky130_a_tran.raw v(in) v(out) avg_pw_total

  dc Vin 0 1 0.00001
  save all
  write tb_inv_sky130_a_DC.raw v(in) v(out)

  exit 0
.endc


**** end user architecture code
**.ends

* expanding   symbol:  inv_sky130_a.sym # of pins=2
** sym_path: /Users/miguelcorrea/Desktop/MA2_project/Amplifier_Inv/xschem/inv_sky130_a.sym
** sch_path: /Users/miguelcorrea/Desktop/MA2_project/Amplifier_Inv/xschem/inv_sky130_a.sch
.subckt inv_sky130_a out in
*.ipin in
*.opin out
x1 test in VCC VSS not W_N=250 L_N=1 W_P=200 L_P=0.25 m=1
XC1 out GND sky130_fd_pr__cap_mim_m3_1 W=55 L=55 MF=5 m=5
XR1 test in GND sky130_fd_pr__res_xhigh_po W=1 L=90 mult=1 m=1
XR2 out test GND sky130_fd_pr__res_xhigh_po W=1 L=50 mult=1 m=1
.ends


* expanding   symbol:  sky130_tests/not.sym # of pins=2
** sym_path: /usr/local/share/pdk/sky130A/libs.tech/xschem/sky130_tests/not.sym
** sch_path: /usr/local/share/pdk/sky130A/libs.tech/xschem/sky130_tests/not.sch
.subckt not y a VCCPIN VSSPIN     W_N=1 L_N=0.15 W_P=2 L_P=0.15
*.opin y
*.ipin a
XM1 y a VSSPIN VSSPIN sky130_fd_pr__nfet_01v8 L=L_N W=W_N nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 y a VCCPIN VCCPIN sky130_fd_pr__pfet_01v8 L=L_P W=W_P nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.GLOBAL VSS
.GLOBAL VCC
.end
