** sch_path: /Users/miguelcorrea/Desktop/MA2_project/Amplifier_Inv/xschem/v4/inv_sky130_a_v4.sch
.subckt inv_sky130_a_v4 VG1 VCC VG2 out in VSS
*.PININFO in:I out:O VG1:I VG2:I VSS:I VCC:I
XC1 in VD1 sky130_fd_pr__cap_mim_m3_1 W=26 L=26 m=1
XM4 VS1 VD1 VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=250 nf=10 m=1
XM5 VS1 VD1 VCC VCC sky130_fd_pr__pfet_01v8 L=0.25 W=200 nf=8 m=1
XM2 VS1 VG2 out VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=1
XM3 VSS out VSS VSS sky130_fd_pr__nfet_01v8 L=10 W=100 nf=4 m=1
XM1 VD1 VG1 VS1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt


**** end user architecture code
.ends
.end
